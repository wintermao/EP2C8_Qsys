// nios2.v

// Generated using ACDS version 13.0 156 at 2018.05.12.09:59:33

`timescale 1 ps / 1 ps
module nios2 (
		input  wire        clk_clk,                  //           clk.clk
		input  wire        reset_reset_n,            //         reset.reset_n
		output wire [11:0] sdram_addr,               //         sdram.addr
		output wire [1:0]  sdram_ba,                 //              .ba
		output wire        sdram_cas_n,              //              .cas_n
		output wire        sdram_cke,                //              .cke
		output wire        sdram_cs_n,               //              .cs_n
		inout  wire [15:0] sdram_dq,                 //              .dq
		output wire [1:0]  sdram_dqm,                //              .dqm
		output wire        sdram_ras_n,              //              .ras_n
		output wire        sdram_we_n,               //              .we_n
		output wire        sdram_clk_clk,            //     sdram_clk.clk
		input  wire        uart1_rxd,                //         uart1.rxd
		output wire        uart1_txd,                //              .txd
		input  wire        uart2_rxd,                //         uart2.rxd
		output wire        uart2_txd,                //              .txd
		input  wire        uart3_rxd,                //         uart3.rxd
		output wire        uart3_txd,                //              .txd
		output wire [4:0]  led_export,               //           led.export
		input  wire [2:0]  key_export,               //           key.export
		inout  wire        oc_i2c_master_scl_pad_io, // oc_i2c_master.scl_pad_io
		inout  wire        oc_i2c_master_sda_pad_io  //              .sda_pad_io
	);

	wire          altpll_c0_clk;                                                                                     // altpll:c0 -> [addr_router:clk, addr_router_001:clk, addr_router_002:clk, addr_router_003:clk, addr_router_004:clk, burst_adapter:clk, burst_adapter_001:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_demux_004:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, cmd_xbar_mux_010:clk, cmd_xbar_mux_015:clk, crosser:in_clk, crosser_001:out_clk, dma_0:clk, dma_0_control_port_slave_translator:clk, dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:clk, dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dma_0_read_master_translator:clk, dma_0_read_master_translator_avalon_universal_master_0_agent:clk, dma_0_write_master_translator:clk, dma_0_write_master_translator_avalon_universal_master_0_agent:clk, epcs_flash:clk, epcs_flash_epcs_control_port_translator:clk, epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:clk, epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, irq_mapper:clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, master_0:clk_clk, master_0_master_translator:clk, master_0_master_translator_avalon_universal_master_0_agent:clk, nios2:clk, nios2_data_master_translator:clk, nios2_data_master_translator_avalon_universal_master_0_agent:clk, nios2_instruction_master_translator:clk, nios2_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_jtag_debug_module_translator:clk, nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, oc_i2c_master_0:wb_clk_i, oc_i2c_master_0_s1_translator:clk, oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:clk, oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_ram:clk, onchip_ram_s1_translator:clk, onchip_ram_s1_translator_avalon_universal_slave_0_agent:clk, onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_key:clk, pio_key_s1_translator:clk, pio_key_s1_translator_avalon_universal_slave_0_agent:clk, pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_led:clk, pio_led_s1_translator:clk, pio_led_s1_translator_avalon_universal_slave_0_agent:clk, pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rsp_xbar_mux_002:clk, rst_controller:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sysid:clock, sysid_control_slave_translator:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, systimer:clk, systimer_s1_translator:clk, systimer_s1_translator_avalon_universal_slave_0_agent:clk, systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timestamp:clk, timestamp_s1_translator:clk, timestamp_s1_translator_avalon_universal_slave_0_agent:clk, timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, uart1:clk, uart1_s1_translator:clk, uart1_s1_translator_avalon_universal_slave_0_agent:clk, uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, uart2:clk, uart2_s1_translator:clk, uart2_s1_translator_avalon_universal_slave_0_agent:clk, uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, uart3:clk, uart3_s1_translator:clk, uart3_s1_translator_avalon_universal_slave_0_agent:clk, uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, width_adapter_008:clk, width_adapter_009:clk, width_adapter_010:clk, width_adapter_011:clk]
	wire          nios2_instruction_master_waitrequest;                                                              // nios2_instruction_master_translator:av_waitrequest -> nios2:i_waitrequest
	wire   [24:0] nios2_instruction_master_address;                                                                  // nios2:i_address -> nios2_instruction_master_translator:av_address
	wire          nios2_instruction_master_read;                                                                     // nios2:i_read -> nios2_instruction_master_translator:av_read
	wire   [31:0] nios2_instruction_master_readdata;                                                                 // nios2_instruction_master_translator:av_readdata -> nios2:i_readdata
	wire          nios2_data_master_waitrequest;                                                                     // nios2_data_master_translator:av_waitrequest -> nios2:d_waitrequest
	wire   [31:0] nios2_data_master_writedata;                                                                       // nios2:d_writedata -> nios2_data_master_translator:av_writedata
	wire   [24:0] nios2_data_master_address;                                                                         // nios2:d_address -> nios2_data_master_translator:av_address
	wire          nios2_data_master_write;                                                                           // nios2:d_write -> nios2_data_master_translator:av_write
	wire          nios2_data_master_read;                                                                            // nios2:d_read -> nios2_data_master_translator:av_read
	wire   [31:0] nios2_data_master_readdata;                                                                        // nios2_data_master_translator:av_readdata -> nios2:d_readdata
	wire          nios2_data_master_debugaccess;                                                                     // nios2:jtag_debug_module_debugaccess_to_roms -> nios2_data_master_translator:av_debugaccess
	wire    [3:0] nios2_data_master_byteenable;                                                                      // nios2:d_byteenable -> nios2_data_master_translator:av_byteenable
	wire          master_0_master_waitrequest;                                                                       // master_0_master_translator:av_waitrequest -> master_0:master_waitrequest
	wire   [31:0] master_0_master_writedata;                                                                         // master_0:master_writedata -> master_0_master_translator:av_writedata
	wire   [31:0] master_0_master_address;                                                                           // master_0:master_address -> master_0_master_translator:av_address
	wire          master_0_master_write;                                                                             // master_0:master_write -> master_0_master_translator:av_write
	wire          master_0_master_read;                                                                              // master_0:master_read -> master_0_master_translator:av_read
	wire   [31:0] master_0_master_readdata;                                                                          // master_0_master_translator:av_readdata -> master_0:master_readdata
	wire    [3:0] master_0_master_byteenable;                                                                        // master_0:master_byteenable -> master_0_master_translator:av_byteenable
	wire          master_0_master_readdatavalid;                                                                     // master_0_master_translator:av_readdatavalid -> master_0:master_readdatavalid
	wire          dma_0_write_master_waitrequest;                                                                    // dma_0_write_master_translator:av_waitrequest -> dma_0:write_waitrequest
	wire   [15:0] dma_0_write_master_writedata;                                                                      // dma_0:write_writedata -> dma_0_write_master_translator:av_writedata
	wire   [24:0] dma_0_write_master_address;                                                                        // dma_0:write_address -> dma_0_write_master_translator:av_address
	wire          dma_0_write_master_chipselect;                                                                     // dma_0:write_chipselect -> dma_0_write_master_translator:av_chipselect
	wire          dma_0_write_master_write;                                                                          // dma_0:write_write_n -> dma_0_write_master_translator:av_write
	wire    [1:0] dma_0_write_master_byteenable;                                                                     // dma_0:write_byteenable -> dma_0_write_master_translator:av_byteenable
	wire          dma_0_read_master_waitrequest;                                                                     // dma_0_read_master_translator:av_waitrequest -> dma_0:read_waitrequest
	wire   [23:0] dma_0_read_master_address;                                                                         // dma_0:read_address -> dma_0_read_master_translator:av_address
	wire          dma_0_read_master_chipselect;                                                                      // dma_0:read_chipselect -> dma_0_read_master_translator:av_chipselect
	wire          dma_0_read_master_read;                                                                            // dma_0:read_read_n -> dma_0_read_master_translator:av_read
	wire   [15:0] dma_0_read_master_readdata;                                                                        // dma_0_read_master_translator:av_readdata -> dma_0:read_readdata
	wire          dma_0_read_master_readdatavalid;                                                                   // dma_0_read_master_translator:av_readdatavalid -> dma_0:read_readdatavalid
	wire          nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                // nios2:jtag_debug_module_waitrequest -> nios2_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                  // nios2_jtag_debug_module_translator:av_writedata -> nios2:jtag_debug_module_writedata
	wire    [8:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_address;                                    // nios2_jtag_debug_module_translator:av_address -> nios2:jtag_debug_module_address
	wire          nios2_jtag_debug_module_translator_avalon_anti_slave_0_write;                                      // nios2_jtag_debug_module_translator:av_write -> nios2:jtag_debug_module_write
	wire          nios2_jtag_debug_module_translator_avalon_anti_slave_0_read;                                       // nios2_jtag_debug_module_translator:av_read -> nios2:jtag_debug_module_read
	wire   [31:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                   // nios2:jtag_debug_module_readdata -> nios2_jtag_debug_module_translator:av_readdata
	wire          nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                // nios2_jtag_debug_module_translator:av_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire    [3:0] nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                 // nios2_jtag_debug_module_translator:av_byteenable -> nios2:jtag_debug_module_byteenable
	wire   [15:0] onchip_ram_s1_translator_avalon_anti_slave_0_writedata;                                            // onchip_ram_s1_translator:av_writedata -> onchip_ram:writedata
	wire   [10:0] onchip_ram_s1_translator_avalon_anti_slave_0_address;                                              // onchip_ram_s1_translator:av_address -> onchip_ram:address
	wire          onchip_ram_s1_translator_avalon_anti_slave_0_chipselect;                                           // onchip_ram_s1_translator:av_chipselect -> onchip_ram:chipselect
	wire          onchip_ram_s1_translator_avalon_anti_slave_0_clken;                                                // onchip_ram_s1_translator:av_clken -> onchip_ram:clken
	wire          onchip_ram_s1_translator_avalon_anti_slave_0_write;                                                // onchip_ram_s1_translator:av_write -> onchip_ram:write
	wire   [15:0] onchip_ram_s1_translator_avalon_anti_slave_0_readdata;                                             // onchip_ram:readdata -> onchip_ram_s1_translator:av_readdata
	wire    [1:0] onchip_ram_s1_translator_avalon_anti_slave_0_byteenable;                                           // onchip_ram_s1_translator:av_byteenable -> onchip_ram:byteenable
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                               // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                 // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [21:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                   // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                     // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                      // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                  // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                             // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire   [31:0] epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_writedata;                             // epcs_flash_epcs_control_port_translator:av_writedata -> epcs_flash:writedata
	wire    [8:0] epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_address;                               // epcs_flash_epcs_control_port_translator:av_address -> epcs_flash:address
	wire          epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_chipselect;                            // epcs_flash_epcs_control_port_translator:av_chipselect -> epcs_flash:chipselect
	wire          epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_write;                                 // epcs_flash_epcs_control_port_translator:av_write -> epcs_flash:write_n
	wire          epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_read;                                  // epcs_flash_epcs_control_port_translator:av_read -> epcs_flash:read_n
	wire   [31:0] epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_readdata;                              // epcs_flash:readdata -> epcs_flash_epcs_control_port_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                        // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                       // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                            // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                              // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                             // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                  // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                   // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                               // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] altpll_pll_slave_translator_avalon_anti_slave_0_writedata;                                         // altpll_pll_slave_translator:av_writedata -> altpll:writedata
	wire    [1:0] altpll_pll_slave_translator_avalon_anti_slave_0_address;                                           // altpll_pll_slave_translator:av_address -> altpll:address
	wire          altpll_pll_slave_translator_avalon_anti_slave_0_write;                                             // altpll_pll_slave_translator:av_write -> altpll:write
	wire          altpll_pll_slave_translator_avalon_anti_slave_0_read;                                              // altpll_pll_slave_translator:av_read -> altpll:read
	wire   [31:0] altpll_pll_slave_translator_avalon_anti_slave_0_readdata;                                          // altpll:readdata -> altpll_pll_slave_translator:av_readdata
	wire   [15:0] systimer_s1_translator_avalon_anti_slave_0_writedata;                                              // systimer_s1_translator:av_writedata -> systimer:writedata
	wire    [2:0] systimer_s1_translator_avalon_anti_slave_0_address;                                                // systimer_s1_translator:av_address -> systimer:address
	wire          systimer_s1_translator_avalon_anti_slave_0_chipselect;                                             // systimer_s1_translator:av_chipselect -> systimer:chipselect
	wire          systimer_s1_translator_avalon_anti_slave_0_write;                                                  // systimer_s1_translator:av_write -> systimer:write_n
	wire   [15:0] systimer_s1_translator_avalon_anti_slave_0_readdata;                                               // systimer:readdata -> systimer_s1_translator:av_readdata
	wire   [15:0] timestamp_s1_translator_avalon_anti_slave_0_writedata;                                             // timestamp_s1_translator:av_writedata -> timestamp:writedata
	wire    [2:0] timestamp_s1_translator_avalon_anti_slave_0_address;                                               // timestamp_s1_translator:av_address -> timestamp:address
	wire          timestamp_s1_translator_avalon_anti_slave_0_chipselect;                                            // timestamp_s1_translator:av_chipselect -> timestamp:chipselect
	wire          timestamp_s1_translator_avalon_anti_slave_0_write;                                                 // timestamp_s1_translator:av_write -> timestamp:write_n
	wire   [15:0] timestamp_s1_translator_avalon_anti_slave_0_readdata;                                              // timestamp:readdata -> timestamp_s1_translator:av_readdata
	wire   [15:0] uart1_s1_translator_avalon_anti_slave_0_writedata;                                                 // uart1_s1_translator:av_writedata -> uart1:writedata
	wire    [2:0] uart1_s1_translator_avalon_anti_slave_0_address;                                                   // uart1_s1_translator:av_address -> uart1:address
	wire          uart1_s1_translator_avalon_anti_slave_0_chipselect;                                                // uart1_s1_translator:av_chipselect -> uart1:chipselect
	wire          uart1_s1_translator_avalon_anti_slave_0_write;                                                     // uart1_s1_translator:av_write -> uart1:write_n
	wire          uart1_s1_translator_avalon_anti_slave_0_read;                                                      // uart1_s1_translator:av_read -> uart1:read_n
	wire   [15:0] uart1_s1_translator_avalon_anti_slave_0_readdata;                                                  // uart1:readdata -> uart1_s1_translator:av_readdata
	wire          uart1_s1_translator_avalon_anti_slave_0_begintransfer;                                             // uart1_s1_translator:av_begintransfer -> uart1:begintransfer
	wire   [15:0] uart2_s1_translator_avalon_anti_slave_0_writedata;                                                 // uart2_s1_translator:av_writedata -> uart2:writedata
	wire    [2:0] uart2_s1_translator_avalon_anti_slave_0_address;                                                   // uart2_s1_translator:av_address -> uart2:address
	wire          uart2_s1_translator_avalon_anti_slave_0_chipselect;                                                // uart2_s1_translator:av_chipselect -> uart2:chipselect
	wire          uart2_s1_translator_avalon_anti_slave_0_write;                                                     // uart2_s1_translator:av_write -> uart2:write_n
	wire          uart2_s1_translator_avalon_anti_slave_0_read;                                                      // uart2_s1_translator:av_read -> uart2:read_n
	wire   [15:0] uart2_s1_translator_avalon_anti_slave_0_readdata;                                                  // uart2:readdata -> uart2_s1_translator:av_readdata
	wire          uart2_s1_translator_avalon_anti_slave_0_begintransfer;                                             // uart2_s1_translator:av_begintransfer -> uart2:begintransfer
	wire   [15:0] uart3_s1_translator_avalon_anti_slave_0_writedata;                                                 // uart3_s1_translator:av_writedata -> uart3:writedata
	wire    [2:0] uart3_s1_translator_avalon_anti_slave_0_address;                                                   // uart3_s1_translator:av_address -> uart3:address
	wire          uart3_s1_translator_avalon_anti_slave_0_chipselect;                                                // uart3_s1_translator:av_chipselect -> uart3:chipselect
	wire          uart3_s1_translator_avalon_anti_slave_0_write;                                                     // uart3_s1_translator:av_write -> uart3:write_n
	wire          uart3_s1_translator_avalon_anti_slave_0_read;                                                      // uart3_s1_translator:av_read -> uart3:read_n
	wire   [15:0] uart3_s1_translator_avalon_anti_slave_0_readdata;                                                  // uart3:readdata -> uart3_s1_translator:av_readdata
	wire          uart3_s1_translator_avalon_anti_slave_0_begintransfer;                                             // uart3_s1_translator:av_begintransfer -> uart3:begintransfer
	wire   [31:0] pio_led_s1_translator_avalon_anti_slave_0_writedata;                                               // pio_led_s1_translator:av_writedata -> pio_led:writedata
	wire    [2:0] pio_led_s1_translator_avalon_anti_slave_0_address;                                                 // pio_led_s1_translator:av_address -> pio_led:address
	wire          pio_led_s1_translator_avalon_anti_slave_0_chipselect;                                              // pio_led_s1_translator:av_chipselect -> pio_led:chipselect
	wire          pio_led_s1_translator_avalon_anti_slave_0_write;                                                   // pio_led_s1_translator:av_write -> pio_led:write_n
	wire   [31:0] pio_led_s1_translator_avalon_anti_slave_0_readdata;                                                // pio_led:readdata -> pio_led_s1_translator:av_readdata
	wire   [31:0] pio_key_s1_translator_avalon_anti_slave_0_writedata;                                               // pio_key_s1_translator:av_writedata -> pio_key:writedata
	wire    [1:0] pio_key_s1_translator_avalon_anti_slave_0_address;                                                 // pio_key_s1_translator:av_address -> pio_key:address
	wire          pio_key_s1_translator_avalon_anti_slave_0_chipselect;                                              // pio_key_s1_translator:av_chipselect -> pio_key:chipselect
	wire          pio_key_s1_translator_avalon_anti_slave_0_write;                                                   // pio_key_s1_translator:av_write -> pio_key:write_n
	wire   [31:0] pio_key_s1_translator_avalon_anti_slave_0_readdata;                                                // pio_key:readdata -> pio_key_s1_translator:av_readdata
	wire          oc_i2c_master_0_s1_translator_avalon_anti_slave_0_waitrequest;                                     // oc_i2c_master_0:wb_ack_o -> oc_i2c_master_0_s1_translator:av_waitrequest
	wire   [31:0] oc_i2c_master_0_s1_translator_avalon_anti_slave_0_writedata;                                       // oc_i2c_master_0_s1_translator:av_writedata -> oc_i2c_master_0:wb_dat_i
	wire    [2:0] oc_i2c_master_0_s1_translator_avalon_anti_slave_0_address;                                         // oc_i2c_master_0_s1_translator:av_address -> oc_i2c_master_0:wb_adr_i
	wire          oc_i2c_master_0_s1_translator_avalon_anti_slave_0_chipselect;                                      // oc_i2c_master_0_s1_translator:av_chipselect -> oc_i2c_master_0:wb_cyc_i
	wire          oc_i2c_master_0_s1_translator_avalon_anti_slave_0_write;                                           // oc_i2c_master_0_s1_translator:av_write -> oc_i2c_master_0:wb_we_i
	wire   [31:0] oc_i2c_master_0_s1_translator_avalon_anti_slave_0_readdata;                                        // oc_i2c_master_0:wb_dat_o -> oc_i2c_master_0_s1_translator:av_readdata
	wire          oc_i2c_master_0_s1_translator_avalon_anti_slave_0_begintransfer;                                   // oc_i2c_master_0_s1_translator:av_begintransfer -> oc_i2c_master_0:wb_stb_i
	wire   [31:0] dma_0_control_port_slave_translator_avalon_anti_slave_0_writedata;                                 // dma_0_control_port_slave_translator:av_writedata -> dma_0:dma_ctl_writedata
	wire    [2:0] dma_0_control_port_slave_translator_avalon_anti_slave_0_address;                                   // dma_0_control_port_slave_translator:av_address -> dma_0:dma_ctl_address
	wire          dma_0_control_port_slave_translator_avalon_anti_slave_0_chipselect;                                // dma_0_control_port_slave_translator:av_chipselect -> dma_0:dma_ctl_chipselect
	wire          dma_0_control_port_slave_translator_avalon_anti_slave_0_write;                                     // dma_0_control_port_slave_translator:av_write -> dma_0:dma_ctl_write_n
	wire   [31:0] dma_0_control_port_slave_translator_avalon_anti_slave_0_readdata;                                  // dma_0:dma_ctl_readdata -> dma_0_control_port_slave_translator:av_readdata
	wire          nios2_instruction_master_translator_avalon_universal_master_0_waitrequest;                         // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_instruction_master_translator_avalon_universal_master_0_burstcount;                          // nios2_instruction_master_translator:uav_burstcount -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_instruction_master_translator_avalon_universal_master_0_writedata;                           // nios2_instruction_master_translator:uav_writedata -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_instruction_master_translator_avalon_universal_master_0_address;                             // nios2_instruction_master_translator:uav_address -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_instruction_master_translator_avalon_universal_master_0_lock;                                // nios2_instruction_master_translator:uav_lock -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_instruction_master_translator_avalon_universal_master_0_write;                               // nios2_instruction_master_translator:uav_write -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_instruction_master_translator_avalon_universal_master_0_read;                                // nios2_instruction_master_translator:uav_read -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_instruction_master_translator_avalon_universal_master_0_readdata;                            // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_instruction_master_translator:uav_readdata
	wire          nios2_instruction_master_translator_avalon_universal_master_0_debugaccess;                         // nios2_instruction_master_translator:uav_debugaccess -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_instruction_master_translator_avalon_universal_master_0_byteenable;                          // nios2_instruction_master_translator:uav_byteenable -> nios2_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid;                       // nios2_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_instruction_master_translator:uav_readdatavalid
	wire          nios2_data_master_translator_avalon_universal_master_0_waitrequest;                                // nios2_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_data_master_translator_avalon_universal_master_0_burstcount;                                 // nios2_data_master_translator:uav_burstcount -> nios2_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_data_master_translator_avalon_universal_master_0_writedata;                                  // nios2_data_master_translator:uav_writedata -> nios2_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_data_master_translator_avalon_universal_master_0_address;                                    // nios2_data_master_translator:uav_address -> nios2_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_data_master_translator_avalon_universal_master_0_lock;                                       // nios2_data_master_translator:uav_lock -> nios2_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_data_master_translator_avalon_universal_master_0_write;                                      // nios2_data_master_translator:uav_write -> nios2_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_data_master_translator_avalon_universal_master_0_read;                                       // nios2_data_master_translator:uav_read -> nios2_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_data_master_translator_avalon_universal_master_0_readdata;                                   // nios2_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_data_master_translator:uav_readdata
	wire          nios2_data_master_translator_avalon_universal_master_0_debugaccess;                                // nios2_data_master_translator:uav_debugaccess -> nios2_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_data_master_translator_avalon_universal_master_0_byteenable;                                 // nios2_data_master_translator:uav_byteenable -> nios2_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_data_master_translator_avalon_universal_master_0_readdatavalid;                              // nios2_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_data_master_translator:uav_readdatavalid
	wire          master_0_master_translator_avalon_universal_master_0_waitrequest;                                  // master_0_master_translator_avalon_universal_master_0_agent:av_waitrequest -> master_0_master_translator:uav_waitrequest
	wire    [2:0] master_0_master_translator_avalon_universal_master_0_burstcount;                                   // master_0_master_translator:uav_burstcount -> master_0_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] master_0_master_translator_avalon_universal_master_0_writedata;                                    // master_0_master_translator:uav_writedata -> master_0_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] master_0_master_translator_avalon_universal_master_0_address;                                      // master_0_master_translator:uav_address -> master_0_master_translator_avalon_universal_master_0_agent:av_address
	wire          master_0_master_translator_avalon_universal_master_0_lock;                                         // master_0_master_translator:uav_lock -> master_0_master_translator_avalon_universal_master_0_agent:av_lock
	wire          master_0_master_translator_avalon_universal_master_0_write;                                        // master_0_master_translator:uav_write -> master_0_master_translator_avalon_universal_master_0_agent:av_write
	wire          master_0_master_translator_avalon_universal_master_0_read;                                         // master_0_master_translator:uav_read -> master_0_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] master_0_master_translator_avalon_universal_master_0_readdata;                                     // master_0_master_translator_avalon_universal_master_0_agent:av_readdata -> master_0_master_translator:uav_readdata
	wire          master_0_master_translator_avalon_universal_master_0_debugaccess;                                  // master_0_master_translator:uav_debugaccess -> master_0_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] master_0_master_translator_avalon_universal_master_0_byteenable;                                   // master_0_master_translator:uav_byteenable -> master_0_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          master_0_master_translator_avalon_universal_master_0_readdatavalid;                                // master_0_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> master_0_master_translator:uav_readdatavalid
	wire          dma_0_read_master_translator_avalon_universal_master_0_waitrequest;                                // dma_0_read_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_0_read_master_translator:uav_waitrequest
	wire    [1:0] dma_0_read_master_translator_avalon_universal_master_0_burstcount;                                 // dma_0_read_master_translator:uav_burstcount -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] dma_0_read_master_translator_avalon_universal_master_0_writedata;                                  // dma_0_read_master_translator:uav_writedata -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] dma_0_read_master_translator_avalon_universal_master_0_address;                                    // dma_0_read_master_translator:uav_address -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_0_read_master_translator_avalon_universal_master_0_lock;                                       // dma_0_read_master_translator:uav_lock -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_0_read_master_translator_avalon_universal_master_0_write;                                      // dma_0_read_master_translator:uav_write -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_0_read_master_translator_avalon_universal_master_0_read;                                       // dma_0_read_master_translator:uav_read -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] dma_0_read_master_translator_avalon_universal_master_0_readdata;                                   // dma_0_read_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_0_read_master_translator:uav_readdata
	wire          dma_0_read_master_translator_avalon_universal_master_0_debugaccess;                                // dma_0_read_master_translator:uav_debugaccess -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] dma_0_read_master_translator_avalon_universal_master_0_byteenable;                                 // dma_0_read_master_translator:uav_byteenable -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_0_read_master_translator_avalon_universal_master_0_readdatavalid;                              // dma_0_read_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_0_read_master_translator:uav_readdatavalid
	wire          dma_0_write_master_translator_avalon_universal_master_0_waitrequest;                               // dma_0_write_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_0_write_master_translator:uav_waitrequest
	wire    [1:0] dma_0_write_master_translator_avalon_universal_master_0_burstcount;                                // dma_0_write_master_translator:uav_burstcount -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] dma_0_write_master_translator_avalon_universal_master_0_writedata;                                 // dma_0_write_master_translator:uav_writedata -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] dma_0_write_master_translator_avalon_universal_master_0_address;                                   // dma_0_write_master_translator:uav_address -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_0_write_master_translator_avalon_universal_master_0_lock;                                      // dma_0_write_master_translator:uav_lock -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_0_write_master_translator_avalon_universal_master_0_write;                                     // dma_0_write_master_translator:uav_write -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_0_write_master_translator_avalon_universal_master_0_read;                                      // dma_0_write_master_translator:uav_read -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] dma_0_write_master_translator_avalon_universal_master_0_readdata;                                  // dma_0_write_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_0_write_master_translator:uav_readdata
	wire          dma_0_write_master_translator_avalon_universal_master_0_debugaccess;                               // dma_0_write_master_translator:uav_debugaccess -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] dma_0_write_master_translator_avalon_universal_master_0_byteenable;                                // dma_0_write_master_translator:uav_byteenable -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_0_write_master_translator_avalon_universal_master_0_readdatavalid;                             // dma_0_write_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_0_write_master_translator:uav_readdatavalid
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                  // nios2_jtag_debug_module_translator:uav_waitrequest -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                   // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                    // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_jtag_debug_module_translator:uav_writedata
	wire   [31:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                      // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_jtag_debug_module_translator:uav_address
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                        // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_jtag_debug_module_translator:uav_write
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                         // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_jtag_debug_module_translator:uav_lock
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                         // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                     // nios2_jtag_debug_module_translator:uav_readdata -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                // nios2_jtag_debug_module_translator:uav_readdatavalid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                  // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                   // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_jtag_debug_module_translator:uav_byteenable
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;           // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                 // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;         // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                  // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                 // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;        // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;              // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;      // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;               // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;              // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;            // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;             // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;            // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // onchip_ram_s1_translator:uav_waitrequest -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_ram_s1_translator:uav_burstcount
	wire   [15:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_ram_s1_translator:uav_writedata
	wire   [31:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_ram_s1_translator:uav_address
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_ram_s1_translator:uav_write
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_ram_s1_translator:uav_lock
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_ram_s1_translator:uav_read
	wire   [15:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // onchip_ram_s1_translator:uav_readdata -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // onchip_ram_s1_translator:uav_readdatavalid -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_ram_s1_translator:uav_debugaccess
	wire    [1:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // onchip_ram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_ram_s1_translator:uav_byteenable
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [89:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [89:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                           // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                            // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                           // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // epcs_flash_epcs_control_port_translator:uav_waitrequest -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount;              // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> epcs_flash_epcs_control_port_translator:uav_burstcount
	wire   [31:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata;               // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> epcs_flash_epcs_control_port_translator:uav_writedata
	wire   [31:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address;                 // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_address -> epcs_flash_epcs_control_port_translator:uav_address
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write;                   // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_write -> epcs_flash_epcs_control_port_translator:uav_write
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock;                    // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> epcs_flash_epcs_control_port_translator:uav_lock
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read;                    // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_read -> epcs_flash_epcs_control_port_translator:uav_read
	wire   [31:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata;                // epcs_flash_epcs_control_port_translator:uav_readdata -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // epcs_flash_epcs_control_port_translator:uav_readdatavalid -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> epcs_flash_epcs_control_port_translator:uav_debugaccess
	wire    [3:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable;              // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> epcs_flash_epcs_control_port_translator:uav_byteenable
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid;            // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data;             // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready;            // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // altpll_pll_slave_translator:uav_waitrequest -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> altpll_pll_slave_translator:uav_burstcount
	wire   [31:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                           // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> altpll_pll_slave_translator:uav_writedata
	wire   [31:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                             // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> altpll_pll_slave_translator:uav_address
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                               // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> altpll_pll_slave_translator:uav_write
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> altpll_pll_slave_translator:uav_lock
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                                // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> altpll_pll_slave_translator:uav_read
	wire   [31:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                            // altpll_pll_slave_translator:uav_readdata -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // altpll_pll_slave_translator:uav_readdatavalid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> altpll_pll_slave_translator:uav_debugaccess
	wire    [3:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // altpll_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> altpll_pll_slave_translator:uav_byteenable
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                         // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                   // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                    // altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                   // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // systimer_s1_translator:uav_waitrequest -> systimer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] systimer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // systimer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> systimer_s1_translator:uav_burstcount
	wire   [31:0] systimer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // systimer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> systimer_s1_translator:uav_writedata
	wire   [31:0] systimer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // systimer_s1_translator_avalon_universal_slave_0_agent:m0_address -> systimer_s1_translator:uav_address
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // systimer_s1_translator_avalon_universal_slave_0_agent:m0_write -> systimer_s1_translator:uav_write
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // systimer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> systimer_s1_translator:uav_lock
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // systimer_s1_translator_avalon_universal_slave_0_agent:m0_read -> systimer_s1_translator:uav_read
	wire   [31:0] systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // systimer_s1_translator:uav_readdata -> systimer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // systimer_s1_translator:uav_readdatavalid -> systimer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // systimer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> systimer_s1_translator:uav_debugaccess
	wire    [3:0] systimer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // systimer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> systimer_s1_translator:uav_byteenable
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // systimer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> systimer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // timestamp_s1_translator:uav_waitrequest -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timestamp_s1_translator:uav_burstcount
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timestamp_s1_translator:uav_writedata
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_address -> timestamp_s1_translator:uav_address
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_write -> timestamp_s1_translator:uav_write
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timestamp_s1_translator:uav_lock
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_read -> timestamp_s1_translator:uav_read
	wire   [31:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // timestamp_s1_translator:uav_readdata -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // timestamp_s1_translator:uav_readdatavalid -> timestamp_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timestamp_s1_translator:uav_debugaccess
	wire    [3:0] timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // timestamp_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timestamp_s1_translator:uav_byteenable
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // timestamp_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // uart1_s1_translator:uav_waitrequest -> uart1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] uart1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // uart1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart1_s1_translator:uav_burstcount
	wire   [31:0] uart1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // uart1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart1_s1_translator:uav_writedata
	wire   [31:0] uart1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // uart1_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart1_s1_translator:uav_address
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // uart1_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart1_s1_translator:uav_write
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // uart1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart1_s1_translator:uav_lock
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // uart1_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart1_s1_translator:uav_read
	wire   [31:0] uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // uart1_s1_translator:uav_readdata -> uart1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // uart1_s1_translator:uav_readdatavalid -> uart1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // uart1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart1_s1_translator:uav_debugaccess
	wire    [3:0] uart1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // uart1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart1_s1_translator:uav_byteenable
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // uart1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // uart1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // uart1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // uart1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // uart1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // uart2_s1_translator:uav_waitrequest -> uart2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] uart2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // uart2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart2_s1_translator:uav_burstcount
	wire   [31:0] uart2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // uart2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart2_s1_translator:uav_writedata
	wire   [31:0] uart2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // uart2_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart2_s1_translator:uav_address
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // uart2_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart2_s1_translator:uav_write
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // uart2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart2_s1_translator:uav_lock
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // uart2_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart2_s1_translator:uav_read
	wire   [31:0] uart2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // uart2_s1_translator:uav_readdata -> uart2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // uart2_s1_translator:uav_readdatavalid -> uart2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // uart2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart2_s1_translator:uav_debugaccess
	wire    [3:0] uart2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // uart2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart2_s1_translator:uav_byteenable
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // uart2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // uart2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // uart2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // uart2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // uart2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // uart2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] uart2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // uart2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // uart2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // uart3_s1_translator:uav_waitrequest -> uart3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] uart3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // uart3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart3_s1_translator:uav_burstcount
	wire   [31:0] uart3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // uart3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart3_s1_translator:uav_writedata
	wire   [31:0] uart3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // uart3_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart3_s1_translator:uav_address
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // uart3_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart3_s1_translator:uav_write
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // uart3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart3_s1_translator:uav_lock
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // uart3_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart3_s1_translator:uav_read
	wire   [31:0] uart3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // uart3_s1_translator:uav_readdata -> uart3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // uart3_s1_translator:uav_readdatavalid -> uart3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // uart3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart3_s1_translator:uav_debugaccess
	wire    [3:0] uart3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // uart3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart3_s1_translator:uav_byteenable
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // uart3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // uart3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // uart3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // uart3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // uart3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // uart3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] uart3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // uart3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // uart3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // pio_led_s1_translator:uav_waitrequest -> pio_led_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_led_s1_translator:uav_burstcount
	wire   [31:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_led_s1_translator:uav_writedata
	wire   [31:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_led_s1_translator:uav_address
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_led_s1_translator:uav_write
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_led_s1_translator:uav_lock
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_led_s1_translator:uav_read
	wire   [31:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // pio_led_s1_translator:uav_readdata -> pio_led_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // pio_led_s1_translator:uav_readdatavalid -> pio_led_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_led_s1_translator:uav_debugaccess
	wire    [3:0] pio_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // pio_led_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_led_s1_translator:uav_byteenable
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // pio_led_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // pio_key_s1_translator:uav_waitrequest -> pio_key_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_key_s1_translator:uav_burstcount
	wire   [31:0] pio_key_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_key_s1_translator:uav_writedata
	wire   [31:0] pio_key_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_key_s1_translator:uav_address
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_key_s1_translator:uav_write
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_key_s1_translator:uav_lock
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_key_s1_translator:uav_read
	wire   [31:0] pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // pio_key_s1_translator:uav_readdata -> pio_key_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // pio_key_s1_translator:uav_readdatavalid -> pio_key_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_key_s1_translator:uav_debugaccess
	wire    [3:0] pio_key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // pio_key_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_key_s1_translator:uav_byteenable
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // pio_key_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // pio_key_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // pio_key_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // pio_key_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_key_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_key_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_key_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // pio_key_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_key_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                       // oc_i2c_master_0_s1_translator:uav_waitrequest -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                        // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> oc_i2c_master_0_s1_translator:uav_burstcount
	wire   [31:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                         // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> oc_i2c_master_0_s1_translator:uav_writedata
	wire   [31:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                           // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> oc_i2c_master_0_s1_translator:uav_address
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                             // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> oc_i2c_master_0_s1_translator:uav_write
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                              // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> oc_i2c_master_0_s1_translator:uav_lock
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                              // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> oc_i2c_master_0_s1_translator:uav_read
	wire   [31:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                          // oc_i2c_master_0_s1_translator:uav_readdata -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                     // oc_i2c_master_0_s1_translator:uav_readdatavalid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                       // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> oc_i2c_master_0_s1_translator:uav_debugaccess
	wire    [3:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                        // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> oc_i2c_master_0_s1_translator:uav_byteenable
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                      // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;              // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                       // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                      // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;             // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                   // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;           // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                    // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                   // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                 // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                  // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                 // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // dma_0_control_port_slave_translator:uav_waitrequest -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> dma_0_control_port_slave_translator:uav_burstcount
	wire   [31:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                   // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> dma_0_control_port_slave_translator:uav_writedata
	wire   [31:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                     // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> dma_0_control_port_slave_translator:uav_address
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                       // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> dma_0_control_port_slave_translator:uav_write
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                        // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> dma_0_control_port_slave_translator:uav_lock
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                        // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> dma_0_control_port_slave_translator:uav_read
	wire   [31:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                    // dma_0_control_port_slave_translator:uav_readdata -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // dma_0_control_port_slave_translator:uav_readdatavalid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dma_0_control_port_slave_translator:uav_debugaccess
	wire    [3:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> dma_0_control_port_slave_translator:uav_byteenable
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                 // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                      // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;              // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [106:0] nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                       // nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                      // addr_router:sink_ready -> nios2_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // nios2_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid;                             // nios2_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // nios2_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [106:0] nios2_data_master_translator_avalon_universal_master_0_agent_cp_data;                              // nios2_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_001:sink_ready -> nios2_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // master_0_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_valid;                               // master_0_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // master_0_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [106:0] master_0_master_translator_avalon_universal_master_0_agent_cp_data;                                // master_0_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router_002:sink_ready -> master_0_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_valid;                             // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire   [88:0] dma_0_read_master_translator_avalon_universal_master_0_agent_cp_data;                              // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_003:sink_ready -> dma_0_read_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_valid;                            // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire   [88:0] dma_0_write_master_translator_avalon_universal_master_0_agent_cp_data;                             // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router_004:sink_ready -> dma_0_write_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                  // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                        // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [106:0] nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                         // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                        // id_router:sink_ready -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [88:0] onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // onchip_ram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_001:sink_ready -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire   [88:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_002:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid;                   // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [106:0] epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data;                    // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [106:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_004:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [106:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_005:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                               // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [106:0] altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                                // altpll_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_006:sink_ready -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // systimer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // systimer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // systimer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [106:0] systimer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // systimer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          systimer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_007:sink_ready -> systimer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [106:0] timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // timestamp_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_008:sink_ready -> timestamp_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // uart1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // uart1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // uart1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [106:0] uart1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // uart1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          uart1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_009:sink_ready -> uart1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // uart2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // uart2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // uart2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [106:0] uart2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // uart2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          uart2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_010:sink_ready -> uart2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // uart3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // uart3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // uart3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [106:0] uart3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // uart3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          uart3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_011:sink_ready -> uart3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [106:0] pio_led_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // pio_led_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          pio_led_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_012:sink_ready -> pio_led_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // pio_key_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // pio_key_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // pio_key_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [106:0] pio_key_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // pio_key_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          pio_key_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_013:sink_ready -> pio_key_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                       // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                             // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                     // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [106:0] oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                              // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                             // id_router_014:sink_ready -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                       // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire  [106:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                        // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_015:sink_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_002_src_endofpacket;                                                                   // addr_router_002:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_002_src_valid;                                                                         // addr_router_002:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_002_src_startofpacket;                                                                 // addr_router_002:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [106:0] addr_router_002_src_data;                                                                          // addr_router_002:src_data -> limiter:cmd_sink_data
	wire   [15:0] addr_router_002_src_channel;                                                                       // addr_router_002:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_002_src_ready;                                                                         // limiter:cmd_sink_ready -> addr_router_002:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                       // limiter:rsp_src_endofpacket -> master_0_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                             // limiter:rsp_src_valid -> master_0_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                     // limiter:rsp_src_startofpacket -> master_0_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_rsp_src_data;                                                                              // limiter:rsp_src_data -> master_0_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] limiter_rsp_src_channel;                                                                           // limiter:rsp_src_channel -> master_0_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                             // master_0_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                 // burst_adapter:source0_endofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                       // burst_adapter:source0_valid -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                               // burst_adapter:source0_startofpacket -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] burst_adapter_source0_data;                                                                        // burst_adapter:source0_data -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                       // onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [15:0] burst_adapter_source0_channel;                                                                     // burst_adapter:source0_channel -> onchip_ram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                             // burst_adapter_001:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                   // burst_adapter_001:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                           // burst_adapter_001:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [88:0] burst_adapter_001_source0_data;                                                                    // burst_adapter_001:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                   // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [15:0] burst_adapter_001_source0_channel;                                                                 // burst_adapter_001:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                    // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, burst_adapter:reset, burst_adapter_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_010:reset, cmd_xbar_mux_015:reset, crosser:in_reset, crosser_001:out_reset, dma_0:system_reset_n, dma_0_control_port_slave_translator:reset, dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:reset, dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_0_read_master_translator:reset, dma_0_read_master_translator_avalon_universal_master_0_agent:reset, dma_0_write_master_translator:reset, dma_0_write_master_translator_avalon_universal_master_0_agent:reset, epcs_flash:reset_n, epcs_flash_epcs_control_port_translator:reset, epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:reset, epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, irq_mapper:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, master_0_master_translator:reset, master_0_master_translator_avalon_universal_master_0_agent:reset, nios2:reset_n, nios2_data_master_translator:reset, nios2_data_master_translator_avalon_universal_master_0_agent:reset, nios2_instruction_master_translator:reset, nios2_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_jtag_debug_module_translator:reset, nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, oc_i2c_master_0:wb_rst_i, oc_i2c_master_0_s1_translator:reset, oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:reset, oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_ram:reset, onchip_ram_s1_translator:reset, onchip_ram_s1_translator_avalon_universal_slave_0_agent:reset, onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_key:reset_n, pio_key_s1_translator:reset, pio_key_s1_translator_avalon_universal_slave_0_agent:reset, pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_led:reset_n, pio_led_s1_translator:reset, pio_led_s1_translator_avalon_universal_slave_0_agent:reset, pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, systimer:reset_n, systimer_s1_translator:reset, systimer_s1_translator_avalon_universal_slave_0_agent:reset, systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timestamp:reset_n, timestamp_s1_translator:reset, timestamp_s1_translator_avalon_universal_slave_0_agent:reset, timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart1:reset_n, uart1_s1_translator:reset, uart1_s1_translator_avalon_universal_slave_0_agent:reset, uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart2:reset_n, uart2_s1_translator:reset, uart2_s1_translator_avalon_universal_slave_0_agent:reset, uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart3:reset_n, uart3_s1_translator:reset, uart3_s1_translator_avalon_universal_slave_0_agent:reset, uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset, width_adapter_010:reset, width_adapter_011:reset]
	wire          nios2_jtag_debug_module_reset_reset;                                                               // nios2:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                                                // rst_controller_001:reset_out -> [altpll:reset, altpll_pll_slave_translator:reset, altpll_pll_slave_translator_avalon_universal_slave_0_agent:reset, altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser:out_reset, crosser_001:in_reset, id_router_006:reset, rsp_xbar_demux_006:reset]
	wire          rst_controller_002_reset_out_reset;                                                                // rst_controller_002:reset_out -> master_0:clk_reset_reset
	wire          cmd_xbar_demux_src0_endofpacket;                                                                   // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                         // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                 // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src0_data;                                                                          // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [15:0] cmd_xbar_demux_src0_channel;                                                                       // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                         // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src3_endofpacket;                                                                   // cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                         // cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                 // cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_src3_data;                                                                          // cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	wire   [15:0] cmd_xbar_demux_src3_channel;                                                                       // cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src3_ready;                                                                         // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                               // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                     // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                             // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src0_data;                                                                      // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src0_channel;                                                                   // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                     // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                               // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                     // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                             // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src3_data;                                                                      // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	wire   [15:0] cmd_xbar_demux_001_src3_channel;                                                                   // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                     // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                               // cmd_xbar_demux_001:src4_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                     // cmd_xbar_demux_001:src4_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                             // cmd_xbar_demux_001:src4_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src4_data;                                                                      // cmd_xbar_demux_001:src4_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src4_channel;                                                                   // cmd_xbar_demux_001:src4_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                               // cmd_xbar_demux_001:src5_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                     // cmd_xbar_demux_001:src5_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                             // cmd_xbar_demux_001:src5_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src5_data;                                                                      // cmd_xbar_demux_001:src5_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src5_channel;                                                                   // cmd_xbar_demux_001:src5_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                               // cmd_xbar_demux_001:src7_endofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                     // cmd_xbar_demux_001:src7_valid -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                             // cmd_xbar_demux_001:src7_startofpacket -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src7_data;                                                                      // cmd_xbar_demux_001:src7_data -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src7_channel;                                                                   // cmd_xbar_demux_001:src7_channel -> systimer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                               // cmd_xbar_demux_001:src8_endofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                     // cmd_xbar_demux_001:src8_valid -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                             // cmd_xbar_demux_001:src8_startofpacket -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src8_data;                                                                      // cmd_xbar_demux_001:src8_data -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src8_channel;                                                                   // cmd_xbar_demux_001:src8_channel -> timestamp_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                               // cmd_xbar_demux_001:src9_endofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                     // cmd_xbar_demux_001:src9_valid -> uart1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                             // cmd_xbar_demux_001:src9_startofpacket -> uart1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src9_data;                                                                      // cmd_xbar_demux_001:src9_data -> uart1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src9_channel;                                                                   // cmd_xbar_demux_001:src9_channel -> uart1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                              // cmd_xbar_demux_001:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                    // cmd_xbar_demux_001:src10_valid -> cmd_xbar_mux_010:sink0_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                            // cmd_xbar_demux_001:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src10_data;                                                                     // cmd_xbar_demux_001:src10_data -> cmd_xbar_mux_010:sink0_data
	wire   [15:0] cmd_xbar_demux_001_src10_channel;                                                                  // cmd_xbar_demux_001:src10_channel -> cmd_xbar_mux_010:sink0_channel
	wire          cmd_xbar_demux_001_src10_ready;                                                                    // cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux_001:src10_ready
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                              // cmd_xbar_demux_001:src11_endofpacket -> uart3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                    // cmd_xbar_demux_001:src11_valid -> uart3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                            // cmd_xbar_demux_001:src11_startofpacket -> uart3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src11_data;                                                                     // cmd_xbar_demux_001:src11_data -> uart3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src11_channel;                                                                  // cmd_xbar_demux_001:src11_channel -> uart3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                              // cmd_xbar_demux_001:src12_endofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                    // cmd_xbar_demux_001:src12_valid -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                            // cmd_xbar_demux_001:src12_startofpacket -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src12_data;                                                                     // cmd_xbar_demux_001:src12_data -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src12_channel;                                                                  // cmd_xbar_demux_001:src12_channel -> pio_led_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                              // cmd_xbar_demux_001:src13_endofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                    // cmd_xbar_demux_001:src13_valid -> pio_key_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                            // cmd_xbar_demux_001:src13_startofpacket -> pio_key_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src13_data;                                                                     // cmd_xbar_demux_001:src13_data -> pio_key_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src13_channel;                                                                  // cmd_xbar_demux_001:src13_channel -> pio_key_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                              // cmd_xbar_demux_001:src14_endofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                    // cmd_xbar_demux_001:src14_valid -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                            // cmd_xbar_demux_001:src14_startofpacket -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src14_data;                                                                     // cmd_xbar_demux_001:src14_data -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_demux_001_src14_channel;                                                                  // cmd_xbar_demux_001:src14_channel -> oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                              // cmd_xbar_demux_001:src15_endofpacket -> cmd_xbar_mux_015:sink0_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                    // cmd_xbar_demux_001:src15_valid -> cmd_xbar_mux_015:sink0_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                            // cmd_xbar_demux_001:src15_startofpacket -> cmd_xbar_mux_015:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src15_data;                                                                     // cmd_xbar_demux_001:src15_data -> cmd_xbar_mux_015:sink0_data
	wire   [15:0] cmd_xbar_demux_001_src15_channel;                                                                  // cmd_xbar_demux_001:src15_channel -> cmd_xbar_mux_015:sink0_channel
	wire          cmd_xbar_demux_001_src15_ready;                                                                    // cmd_xbar_mux_015:sink0_ready -> cmd_xbar_demux_001:src15_ready
	wire          cmd_xbar_demux_002_src2_endofpacket;                                                               // cmd_xbar_demux_002:src2_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire          cmd_xbar_demux_002_src2_valid;                                                                     // cmd_xbar_demux_002:src2_valid -> cmd_xbar_mux_010:sink1_valid
	wire          cmd_xbar_demux_002_src2_startofpacket;                                                             // cmd_xbar_demux_002:src2_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src2_data;                                                                      // cmd_xbar_demux_002:src2_data -> cmd_xbar_mux_010:sink1_data
	wire   [15:0] cmd_xbar_demux_002_src2_channel;                                                                   // cmd_xbar_demux_002:src2_channel -> cmd_xbar_mux_010:sink1_channel
	wire          cmd_xbar_demux_002_src2_ready;                                                                     // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_002:src2_ready
	wire          cmd_xbar_demux_002_src3_endofpacket;                                                               // cmd_xbar_demux_002:src3_endofpacket -> cmd_xbar_mux_015:sink1_endofpacket
	wire          cmd_xbar_demux_002_src3_valid;                                                                     // cmd_xbar_demux_002:src3_valid -> cmd_xbar_mux_015:sink1_valid
	wire          cmd_xbar_demux_002_src3_startofpacket;                                                             // cmd_xbar_demux_002:src3_startofpacket -> cmd_xbar_mux_015:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src3_data;                                                                      // cmd_xbar_demux_002:src3_data -> cmd_xbar_mux_015:sink1_data
	wire   [15:0] cmd_xbar_demux_002_src3_channel;                                                                   // cmd_xbar_demux_002:src3_channel -> cmd_xbar_mux_015:sink1_channel
	wire          cmd_xbar_demux_002_src3_ready;                                                                     // cmd_xbar_mux_015:sink1_ready -> cmd_xbar_demux_002:src3_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                               // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_002:sink3_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                     // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_002:sink3_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                             // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_002:sink3_startofpacket
	wire   [88:0] cmd_xbar_demux_003_src0_data;                                                                      // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_002:sink3_data
	wire   [15:0] cmd_xbar_demux_003_src0_channel;                                                                   // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_002:sink3_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                     // cmd_xbar_mux_002:sink3_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                               // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_001:sink3_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                     // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_001:sink3_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                             // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_001:sink3_startofpacket
	wire   [88:0] cmd_xbar_demux_004_src0_data;                                                                      // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_001:sink3_data
	wire   [15:0] cmd_xbar_demux_004_src0_channel;                                                                   // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_001:sink3_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                     // cmd_xbar_mux_001:sink3_ready -> cmd_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                   // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                         // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                 // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src0_data;                                                                          // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [15:0] rsp_xbar_demux_src0_channel;                                                                       // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                         // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                   // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                         // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                 // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_src1_data;                                                                          // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [15:0] rsp_xbar_demux_src1_channel;                                                                       // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                         // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src3_endofpacket;                                                               // rsp_xbar_demux_001:src3_endofpacket -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_001_src3_valid;                                                                     // rsp_xbar_demux_001:src3_valid -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_001_src3_startofpacket;                                                             // rsp_xbar_demux_001:src3_startofpacket -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src3_data;                                                                      // rsp_xbar_demux_001:src3_data -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_demux_001_src3_channel;                                                                   // rsp_xbar_demux_001:src3_channel -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_002_src3_endofpacket;                                                               // rsp_xbar_demux_002:src3_endofpacket -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_002_src3_valid;                                                                     // rsp_xbar_demux_002:src3_valid -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_002_src3_startofpacket;                                                             // rsp_xbar_demux_002:src3_startofpacket -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [88:0] rsp_xbar_demux_002_src3_data;                                                                      // rsp_xbar_demux_002:src3_data -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_demux_002_src3_channel;                                                                   // rsp_xbar_demux_002:src3_channel -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                               // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                     // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                             // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src0_data;                                                                      // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire   [15:0] rsp_xbar_demux_003_src0_channel;                                                                   // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                     // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                               // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                     // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                             // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_003_src1_data;                                                                      // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	wire   [15:0] rsp_xbar_demux_003_src1_channel;                                                                   // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                     // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                               // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                     // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                             // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src0_data;                                                                      // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire   [15:0] rsp_xbar_demux_004_src0_channel;                                                                   // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                     // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                               // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                     // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                             // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_005_src0_data;                                                                      // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire   [15:0] rsp_xbar_demux_005_src0_channel;                                                                   // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                     // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                               // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                     // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                             // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [106:0] rsp_xbar_demux_007_src0_data;                                                                      // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire   [15:0] rsp_xbar_demux_007_src0_channel;                                                                   // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                     // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                               // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                     // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                             // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [106:0] rsp_xbar_demux_008_src0_data;                                                                      // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire   [15:0] rsp_xbar_demux_008_src0_channel;                                                                   // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                     // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                               // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                     // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                             // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [106:0] rsp_xbar_demux_009_src0_data;                                                                      // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire   [15:0] rsp_xbar_demux_009_src0_channel;                                                                   // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                     // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                               // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                     // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                             // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [106:0] rsp_xbar_demux_010_src0_data;                                                                      // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire   [15:0] rsp_xbar_demux_010_src0_channel;                                                                   // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                     // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_010_src1_endofpacket;                                                               // rsp_xbar_demux_010:src1_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire          rsp_xbar_demux_010_src1_valid;                                                                     // rsp_xbar_demux_010:src1_valid -> rsp_xbar_mux_002:sink2_valid
	wire          rsp_xbar_demux_010_src1_startofpacket;                                                             // rsp_xbar_demux_010:src1_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_010_src1_data;                                                                      // rsp_xbar_demux_010:src1_data -> rsp_xbar_mux_002:sink2_data
	wire   [15:0] rsp_xbar_demux_010_src1_channel;                                                                   // rsp_xbar_demux_010:src1_channel -> rsp_xbar_mux_002:sink2_channel
	wire          rsp_xbar_demux_010_src1_ready;                                                                     // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_010:src1_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                               // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                     // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                             // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [106:0] rsp_xbar_demux_011_src0_data;                                                                      // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire   [15:0] rsp_xbar_demux_011_src0_channel;                                                                   // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                     // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                               // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                     // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                             // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [106:0] rsp_xbar_demux_012_src0_data;                                                                      // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire   [15:0] rsp_xbar_demux_012_src0_channel;                                                                   // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                     // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                               // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                     // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                             // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [106:0] rsp_xbar_demux_013_src0_data;                                                                      // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire   [15:0] rsp_xbar_demux_013_src0_channel;                                                                   // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                     // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                               // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                     // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                             // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [106:0] rsp_xbar_demux_014_src0_data;                                                                      // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	wire   [15:0] rsp_xbar_demux_014_src0_channel;                                                                   // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                     // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                               // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                     // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                             // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [106:0] rsp_xbar_demux_015_src0_data;                                                                      // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	wire   [15:0] rsp_xbar_demux_015_src0_channel;                                                                   // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                     // rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_015_src1_endofpacket;                                                               // rsp_xbar_demux_015:src1_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire          rsp_xbar_demux_015_src1_valid;                                                                     // rsp_xbar_demux_015:src1_valid -> rsp_xbar_mux_002:sink3_valid
	wire          rsp_xbar_demux_015_src1_startofpacket;                                                             // rsp_xbar_demux_015:src1_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_015_src1_data;                                                                      // rsp_xbar_demux_015:src1_data -> rsp_xbar_mux_002:sink3_data
	wire   [15:0] rsp_xbar_demux_015_src1_channel;                                                                   // rsp_xbar_demux_015:src1_channel -> rsp_xbar_mux_002:sink3_channel
	wire          rsp_xbar_demux_015_src1_ready;                                                                     // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_015:src1_ready
	wire          addr_router_src_endofpacket;                                                                       // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                                             // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                                     // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [106:0] addr_router_src_data;                                                                              // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire   [15:0] addr_router_src_channel;                                                                           // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                                             // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                      // rsp_xbar_mux:src_endofpacket -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                            // rsp_xbar_mux:src_valid -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                    // rsp_xbar_mux:src_startofpacket -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_src_data;                                                                             // rsp_xbar_mux:src_data -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_mux_src_channel;                                                                          // rsp_xbar_mux:src_channel -> nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_src_ready;                                                                            // nios2_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	wire          addr_router_001_src_endofpacket;                                                                   // addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          addr_router_001_src_valid;                                                                         // addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	wire          addr_router_001_src_startofpacket;                                                                 // addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [106:0] addr_router_001_src_data;                                                                          // addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	wire   [15:0] addr_router_001_src_channel;                                                                       // addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	wire          addr_router_001_src_ready;                                                                         // cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                  // rsp_xbar_mux_001:src_endofpacket -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                        // rsp_xbar_mux_001:src_valid -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                // rsp_xbar_mux_001:src_startofpacket -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] rsp_xbar_mux_001_src_data;                                                                         // rsp_xbar_mux_001:src_data -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [15:0] rsp_xbar_mux_001_src_channel;                                                                      // rsp_xbar_mux_001:src_channel -> nios2_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                        // nios2_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	wire          limiter_cmd_src_endofpacket;                                                                       // limiter:cmd_src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                     // limiter:cmd_src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [106:0] limiter_cmd_src_data;                                                                              // limiter:cmd_src_data -> cmd_xbar_demux_002:sink_data
	wire   [15:0] limiter_cmd_src_channel;                                                                           // limiter:cmd_src_channel -> cmd_xbar_demux_002:sink_channel
	wire          limiter_cmd_src_ready;                                                                             // cmd_xbar_demux_002:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                  // rsp_xbar_mux_002:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                        // rsp_xbar_mux_002:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                                // rsp_xbar_mux_002:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_002_src_data;                                                                         // rsp_xbar_mux_002:src_data -> limiter:rsp_sink_data
	wire   [15:0] rsp_xbar_mux_002_src_channel;                                                                      // rsp_xbar_mux_002:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                        // limiter:rsp_sink_ready -> rsp_xbar_mux_002:src_ready
	wire          addr_router_003_src_endofpacket;                                                                   // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                         // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                 // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire   [88:0] addr_router_003_src_data;                                                                          // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire   [15:0] addr_router_003_src_channel;                                                                       // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                         // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_demux_002_src3_ready;                                                                     // dma_0_read_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_002:src3_ready
	wire          addr_router_004_src_endofpacket;                                                                   // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                         // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                 // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire   [88:0] addr_router_004_src_data;                                                                          // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire   [15:0] addr_router_004_src_channel;                                                                       // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                         // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          rsp_xbar_demux_001_src3_ready;                                                                     // dma_0_write_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_001:src3_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                      // cmd_xbar_mux:src_endofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                            // cmd_xbar_mux:src_valid -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                    // cmd_xbar_mux:src_startofpacket -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_src_data;                                                                             // cmd_xbar_mux:src_data -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_src_channel;                                                                          // cmd_xbar_mux:src_channel -> nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                            // nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                         // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                               // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                       // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [106:0] id_router_src_data;                                                                                // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [15:0] id_router_src_channel;                                                                             // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                               // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                  // cmd_xbar_mux_001:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                        // cmd_xbar_mux_001:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                // cmd_xbar_mux_001:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [88:0] cmd_xbar_mux_001_src_data;                                                                         // cmd_xbar_mux_001:src_data -> burst_adapter:sink0_data
	wire   [15:0] cmd_xbar_mux_001_src_channel;                                                                      // cmd_xbar_mux_001:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                        // burst_adapter:sink0_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                     // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                           // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                   // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [88:0] id_router_001_src_data;                                                                            // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [15:0] id_router_001_src_channel;                                                                         // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                           // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                  // cmd_xbar_mux_002:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                        // cmd_xbar_mux_002:src_valid -> burst_adapter_001:sink0_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                // cmd_xbar_mux_002:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [88:0] cmd_xbar_mux_002_src_data;                                                                         // cmd_xbar_mux_002:src_data -> burst_adapter_001:sink0_data
	wire   [15:0] cmd_xbar_mux_002_src_channel;                                                                      // cmd_xbar_mux_002:src_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                        // burst_adapter_001:sink0_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                     // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                           // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                   // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire   [88:0] id_router_002_src_data;                                                                            // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [15:0] id_router_002_src_channel;                                                                         // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                           // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                  // cmd_xbar_mux_003:src_endofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                        // cmd_xbar_mux_003:src_valid -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                // cmd_xbar_mux_003:src_startofpacket -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_003_src_data;                                                                         // cmd_xbar_mux_003:src_data -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_003_src_channel;                                                                      // cmd_xbar_mux_003:src_channel -> epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                        // epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                     // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                           // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                   // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [106:0] id_router_003_src_data;                                                                            // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [15:0] id_router_003_src_channel;                                                                         // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                           // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_001_src4_ready;                                                                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire          id_router_004_src_endofpacket;                                                                     // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                           // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                   // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [106:0] id_router_004_src_data;                                                                            // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [15:0] id_router_004_src_channel;                                                                         // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                           // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_demux_001_src5_ready;                                                                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire          id_router_005_src_endofpacket;                                                                     // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                           // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                   // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [106:0] id_router_005_src_data;                                                                            // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [15:0] id_router_005_src_channel;                                                                         // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                           // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          crosser_out_ready;                                                                                 // altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser:out_ready
	wire          id_router_006_src_endofpacket;                                                                     // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                           // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                   // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [106:0] id_router_006_src_data;                                                                            // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [15:0] id_router_006_src_channel;                                                                         // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                           // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_001_src7_ready;                                                                     // systimer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire          id_router_007_src_endofpacket;                                                                     // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                           // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                   // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [106:0] id_router_007_src_data;                                                                            // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [15:0] id_router_007_src_channel;                                                                         // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                           // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_001_src8_ready;                                                                     // timestamp_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire          id_router_008_src_endofpacket;                                                                     // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                           // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                   // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [106:0] id_router_008_src_data;                                                                            // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [15:0] id_router_008_src_channel;                                                                         // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                           // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_001_src9_ready;                                                                     // uart1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire          id_router_009_src_endofpacket;                                                                     // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                           // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                   // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [106:0] id_router_009_src_data;                                                                            // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [15:0] id_router_009_src_channel;                                                                         // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                           // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_mux_010_src_endofpacket;                                                                  // cmd_xbar_mux_010:src_endofpacket -> uart2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_010_src_valid;                                                                        // cmd_xbar_mux_010:src_valid -> uart2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_010_src_startofpacket;                                                                // cmd_xbar_mux_010:src_startofpacket -> uart2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_010_src_data;                                                                         // cmd_xbar_mux_010:src_data -> uart2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_010_src_channel;                                                                      // cmd_xbar_mux_010:src_channel -> uart2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_010_src_ready;                                                                        // uart2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	wire          id_router_010_src_endofpacket;                                                                     // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                           // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                   // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [106:0] id_router_010_src_data;                                                                            // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [15:0] id_router_010_src_channel;                                                                         // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                           // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_001_src11_ready;                                                                    // uart3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire          id_router_011_src_endofpacket;                                                                     // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                           // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                   // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [106:0] id_router_011_src_data;                                                                            // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [15:0] id_router_011_src_channel;                                                                         // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                           // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_demux_001_src12_ready;                                                                    // pio_led_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire          id_router_012_src_endofpacket;                                                                     // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                           // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                   // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [106:0] id_router_012_src_data;                                                                            // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [15:0] id_router_012_src_channel;                                                                         // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                           // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_demux_001_src13_ready;                                                                    // pio_key_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire          id_router_013_src_endofpacket;                                                                     // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                           // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                   // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [106:0] id_router_013_src_data;                                                                            // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [15:0] id_router_013_src_channel;                                                                         // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                           // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_001_src14_ready;                                                                    // oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	wire          id_router_014_src_endofpacket;                                                                     // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                           // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                   // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [106:0] id_router_014_src_data;                                                                            // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [15:0] id_router_014_src_channel;                                                                         // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                           // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_mux_015_src_endofpacket;                                                                  // cmd_xbar_mux_015:src_endofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_015_src_valid;                                                                        // cmd_xbar_mux_015:src_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_015_src_startofpacket;                                                                // cmd_xbar_mux_015:src_startofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_015_src_data;                                                                         // cmd_xbar_mux_015:src_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] cmd_xbar_mux_015_src_channel;                                                                      // cmd_xbar_mux_015:src_channel -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_015_src_ready;                                                                        // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_015:src_ready
	wire          id_router_015_src_endofpacket;                                                                     // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                           // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                   // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire  [106:0] id_router_015_src_data;                                                                            // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [15:0] id_router_015_src_channel;                                                                         // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                           // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                   // cmd_xbar_demux:src1_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                         // cmd_xbar_demux:src1_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                 // cmd_xbar_demux:src1_startofpacket -> width_adapter:in_startofpacket
	wire  [106:0] cmd_xbar_demux_src1_data;                                                                          // cmd_xbar_demux:src1_data -> width_adapter:in_data
	wire   [15:0] cmd_xbar_demux_src1_channel;                                                                       // cmd_xbar_demux:src1_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src1_ready;                                                                         // width_adapter:in_ready -> cmd_xbar_demux:src1_ready
	wire          width_adapter_src_endofpacket;                                                                     // width_adapter:out_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                           // width_adapter:out_valid -> cmd_xbar_mux_001:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                   // width_adapter:out_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire   [88:0] width_adapter_src_data;                                                                            // width_adapter:out_data -> cmd_xbar_mux_001:sink0_data
	wire          width_adapter_src_ready;                                                                           // cmd_xbar_mux_001:sink0_ready -> width_adapter:out_ready
	wire   [15:0] width_adapter_src_channel;                                                                         // width_adapter:out_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src2_endofpacket;                                                                   // cmd_xbar_demux:src2_endofpacket -> width_adapter_001:in_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                         // cmd_xbar_demux:src2_valid -> width_adapter_001:in_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                 // cmd_xbar_demux:src2_startofpacket -> width_adapter_001:in_startofpacket
	wire  [106:0] cmd_xbar_demux_src2_data;                                                                          // cmd_xbar_demux:src2_data -> width_adapter_001:in_data
	wire   [15:0] cmd_xbar_demux_src2_channel;                                                                       // cmd_xbar_demux:src2_channel -> width_adapter_001:in_channel
	wire          cmd_xbar_demux_src2_ready;                                                                         // width_adapter_001:in_ready -> cmd_xbar_demux:src2_ready
	wire          width_adapter_001_src_endofpacket;                                                                 // width_adapter_001:out_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          width_adapter_001_src_valid;                                                                       // width_adapter_001:out_valid -> cmd_xbar_mux_002:sink0_valid
	wire          width_adapter_001_src_startofpacket;                                                               // width_adapter_001:out_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire   [88:0] width_adapter_001_src_data;                                                                        // width_adapter_001:out_data -> cmd_xbar_mux_002:sink0_data
	wire          width_adapter_001_src_ready;                                                                       // cmd_xbar_mux_002:sink0_ready -> width_adapter_001:out_ready
	wire   [15:0] width_adapter_001_src_channel;                                                                     // width_adapter_001:out_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                               // cmd_xbar_demux_001:src1_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                     // cmd_xbar_demux_001:src1_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                             // cmd_xbar_demux_001:src1_startofpacket -> width_adapter_002:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src1_data;                                                                      // cmd_xbar_demux_001:src1_data -> width_adapter_002:in_data
	wire   [15:0] cmd_xbar_demux_001_src1_channel;                                                                   // cmd_xbar_demux_001:src1_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                     // width_adapter_002:in_ready -> cmd_xbar_demux_001:src1_ready
	wire          width_adapter_002_src_endofpacket;                                                                 // width_adapter_002:out_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          width_adapter_002_src_valid;                                                                       // width_adapter_002:out_valid -> cmd_xbar_mux_001:sink1_valid
	wire          width_adapter_002_src_startofpacket;                                                               // width_adapter_002:out_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire   [88:0] width_adapter_002_src_data;                                                                        // width_adapter_002:out_data -> cmd_xbar_mux_001:sink1_data
	wire          width_adapter_002_src_ready;                                                                       // cmd_xbar_mux_001:sink1_ready -> width_adapter_002:out_ready
	wire   [15:0] width_adapter_002_src_channel;                                                                     // width_adapter_002:out_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                               // cmd_xbar_demux_001:src2_endofpacket -> width_adapter_003:in_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                     // cmd_xbar_demux_001:src2_valid -> width_adapter_003:in_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                             // cmd_xbar_demux_001:src2_startofpacket -> width_adapter_003:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src2_data;                                                                      // cmd_xbar_demux_001:src2_data -> width_adapter_003:in_data
	wire   [15:0] cmd_xbar_demux_001_src2_channel;                                                                   // cmd_xbar_demux_001:src2_channel -> width_adapter_003:in_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                     // width_adapter_003:in_ready -> cmd_xbar_demux_001:src2_ready
	wire          width_adapter_003_src_endofpacket;                                                                 // width_adapter_003:out_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          width_adapter_003_src_valid;                                                                       // width_adapter_003:out_valid -> cmd_xbar_mux_002:sink1_valid
	wire          width_adapter_003_src_startofpacket;                                                               // width_adapter_003:out_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire   [88:0] width_adapter_003_src_data;                                                                        // width_adapter_003:out_data -> cmd_xbar_mux_002:sink1_data
	wire          width_adapter_003_src_ready;                                                                       // cmd_xbar_mux_002:sink1_ready -> width_adapter_003:out_ready
	wire   [15:0] width_adapter_003_src_channel;                                                                     // width_adapter_003:out_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                               // cmd_xbar_demux_002:src0_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                     // cmd_xbar_demux_002:src0_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                             // cmd_xbar_demux_002:src0_startofpacket -> width_adapter_004:in_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src0_data;                                                                      // cmd_xbar_demux_002:src0_data -> width_adapter_004:in_data
	wire   [15:0] cmd_xbar_demux_002_src0_channel;                                                                   // cmd_xbar_demux_002:src0_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                     // width_adapter_004:in_ready -> cmd_xbar_demux_002:src0_ready
	wire          width_adapter_004_src_endofpacket;                                                                 // width_adapter_004:out_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire          width_adapter_004_src_valid;                                                                       // width_adapter_004:out_valid -> cmd_xbar_mux_001:sink2_valid
	wire          width_adapter_004_src_startofpacket;                                                               // width_adapter_004:out_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire   [88:0] width_adapter_004_src_data;                                                                        // width_adapter_004:out_data -> cmd_xbar_mux_001:sink2_data
	wire          width_adapter_004_src_ready;                                                                       // cmd_xbar_mux_001:sink2_ready -> width_adapter_004:out_ready
	wire   [15:0] width_adapter_004_src_channel;                                                                     // width_adapter_004:out_channel -> cmd_xbar_mux_001:sink2_channel
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                               // cmd_xbar_demux_002:src1_endofpacket -> width_adapter_005:in_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                     // cmd_xbar_demux_002:src1_valid -> width_adapter_005:in_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                             // cmd_xbar_demux_002:src1_startofpacket -> width_adapter_005:in_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src1_data;                                                                      // cmd_xbar_demux_002:src1_data -> width_adapter_005:in_data
	wire   [15:0] cmd_xbar_demux_002_src1_channel;                                                                   // cmd_xbar_demux_002:src1_channel -> width_adapter_005:in_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                     // width_adapter_005:in_ready -> cmd_xbar_demux_002:src1_ready
	wire          width_adapter_005_src_endofpacket;                                                                 // width_adapter_005:out_endofpacket -> cmd_xbar_mux_002:sink2_endofpacket
	wire          width_adapter_005_src_valid;                                                                       // width_adapter_005:out_valid -> cmd_xbar_mux_002:sink2_valid
	wire          width_adapter_005_src_startofpacket;                                                               // width_adapter_005:out_startofpacket -> cmd_xbar_mux_002:sink2_startofpacket
	wire   [88:0] width_adapter_005_src_data;                                                                        // width_adapter_005:out_data -> cmd_xbar_mux_002:sink2_data
	wire          width_adapter_005_src_ready;                                                                       // cmd_xbar_mux_002:sink2_ready -> width_adapter_005:out_ready
	wire   [15:0] width_adapter_005_src_channel;                                                                     // width_adapter_005:out_channel -> cmd_xbar_mux_002:sink2_channel
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                               // rsp_xbar_demux_001:src0_endofpacket -> width_adapter_006:in_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                     // rsp_xbar_demux_001:src0_valid -> width_adapter_006:in_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                             // rsp_xbar_demux_001:src0_startofpacket -> width_adapter_006:in_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src0_data;                                                                      // rsp_xbar_demux_001:src0_data -> width_adapter_006:in_data
	wire   [15:0] rsp_xbar_demux_001_src0_channel;                                                                   // rsp_xbar_demux_001:src0_channel -> width_adapter_006:in_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                     // width_adapter_006:in_ready -> rsp_xbar_demux_001:src0_ready
	wire          width_adapter_006_src_endofpacket;                                                                 // width_adapter_006:out_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          width_adapter_006_src_valid;                                                                       // width_adapter_006:out_valid -> rsp_xbar_mux:sink1_valid
	wire          width_adapter_006_src_startofpacket;                                                               // width_adapter_006:out_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [106:0] width_adapter_006_src_data;                                                                        // width_adapter_006:out_data -> rsp_xbar_mux:sink1_data
	wire          width_adapter_006_src_ready;                                                                       // rsp_xbar_mux:sink1_ready -> width_adapter_006:out_ready
	wire   [15:0] width_adapter_006_src_channel;                                                                     // width_adapter_006:out_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                               // rsp_xbar_demux_001:src1_endofpacket -> width_adapter_007:in_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                     // rsp_xbar_demux_001:src1_valid -> width_adapter_007:in_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                             // rsp_xbar_demux_001:src1_startofpacket -> width_adapter_007:in_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src1_data;                                                                      // rsp_xbar_demux_001:src1_data -> width_adapter_007:in_data
	wire   [15:0] rsp_xbar_demux_001_src1_channel;                                                                   // rsp_xbar_demux_001:src1_channel -> width_adapter_007:in_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                     // width_adapter_007:in_ready -> rsp_xbar_demux_001:src1_ready
	wire          width_adapter_007_src_endofpacket;                                                                 // width_adapter_007:out_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          width_adapter_007_src_valid;                                                                       // width_adapter_007:out_valid -> rsp_xbar_mux_001:sink1_valid
	wire          width_adapter_007_src_startofpacket;                                                               // width_adapter_007:out_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [106:0] width_adapter_007_src_data;                                                                        // width_adapter_007:out_data -> rsp_xbar_mux_001:sink1_data
	wire          width_adapter_007_src_ready;                                                                       // rsp_xbar_mux_001:sink1_ready -> width_adapter_007:out_ready
	wire   [15:0] width_adapter_007_src_channel;                                                                     // width_adapter_007:out_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_001_src2_endofpacket;                                                               // rsp_xbar_demux_001:src2_endofpacket -> width_adapter_008:in_endofpacket
	wire          rsp_xbar_demux_001_src2_valid;                                                                     // rsp_xbar_demux_001:src2_valid -> width_adapter_008:in_valid
	wire          rsp_xbar_demux_001_src2_startofpacket;                                                             // rsp_xbar_demux_001:src2_startofpacket -> width_adapter_008:in_startofpacket
	wire   [88:0] rsp_xbar_demux_001_src2_data;                                                                      // rsp_xbar_demux_001:src2_data -> width_adapter_008:in_data
	wire   [15:0] rsp_xbar_demux_001_src2_channel;                                                                   // rsp_xbar_demux_001:src2_channel -> width_adapter_008:in_channel
	wire          rsp_xbar_demux_001_src2_ready;                                                                     // width_adapter_008:in_ready -> rsp_xbar_demux_001:src2_ready
	wire          width_adapter_008_src_endofpacket;                                                                 // width_adapter_008:out_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          width_adapter_008_src_valid;                                                                       // width_adapter_008:out_valid -> rsp_xbar_mux_002:sink0_valid
	wire          width_adapter_008_src_startofpacket;                                                               // width_adapter_008:out_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [106:0] width_adapter_008_src_data;                                                                        // width_adapter_008:out_data -> rsp_xbar_mux_002:sink0_data
	wire          width_adapter_008_src_ready;                                                                       // rsp_xbar_mux_002:sink0_ready -> width_adapter_008:out_ready
	wire   [15:0] width_adapter_008_src_channel;                                                                     // width_adapter_008:out_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                               // rsp_xbar_demux_002:src0_endofpacket -> width_adapter_009:in_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                     // rsp_xbar_demux_002:src0_valid -> width_adapter_009:in_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                             // rsp_xbar_demux_002:src0_startofpacket -> width_adapter_009:in_startofpacket
	wire   [88:0] rsp_xbar_demux_002_src0_data;                                                                      // rsp_xbar_demux_002:src0_data -> width_adapter_009:in_data
	wire   [15:0] rsp_xbar_demux_002_src0_channel;                                                                   // rsp_xbar_demux_002:src0_channel -> width_adapter_009:in_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                     // width_adapter_009:in_ready -> rsp_xbar_demux_002:src0_ready
	wire          width_adapter_009_src_endofpacket;                                                                 // width_adapter_009:out_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          width_adapter_009_src_valid;                                                                       // width_adapter_009:out_valid -> rsp_xbar_mux:sink2_valid
	wire          width_adapter_009_src_startofpacket;                                                               // width_adapter_009:out_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [106:0] width_adapter_009_src_data;                                                                        // width_adapter_009:out_data -> rsp_xbar_mux:sink2_data
	wire          width_adapter_009_src_ready;                                                                       // rsp_xbar_mux:sink2_ready -> width_adapter_009:out_ready
	wire   [15:0] width_adapter_009_src_channel;                                                                     // width_adapter_009:out_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                               // rsp_xbar_demux_002:src1_endofpacket -> width_adapter_010:in_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                     // rsp_xbar_demux_002:src1_valid -> width_adapter_010:in_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                             // rsp_xbar_demux_002:src1_startofpacket -> width_adapter_010:in_startofpacket
	wire   [88:0] rsp_xbar_demux_002_src1_data;                                                                      // rsp_xbar_demux_002:src1_data -> width_adapter_010:in_data
	wire   [15:0] rsp_xbar_demux_002_src1_channel;                                                                   // rsp_xbar_demux_002:src1_channel -> width_adapter_010:in_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                     // width_adapter_010:in_ready -> rsp_xbar_demux_002:src1_ready
	wire          width_adapter_010_src_endofpacket;                                                                 // width_adapter_010:out_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          width_adapter_010_src_valid;                                                                       // width_adapter_010:out_valid -> rsp_xbar_mux_001:sink2_valid
	wire          width_adapter_010_src_startofpacket;                                                               // width_adapter_010:out_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [106:0] width_adapter_010_src_data;                                                                        // width_adapter_010:out_data -> rsp_xbar_mux_001:sink2_data
	wire          width_adapter_010_src_ready;                                                                       // rsp_xbar_mux_001:sink2_ready -> width_adapter_010:out_ready
	wire   [15:0] width_adapter_010_src_channel;                                                                     // width_adapter_010:out_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src2_endofpacket;                                                               // rsp_xbar_demux_002:src2_endofpacket -> width_adapter_011:in_endofpacket
	wire          rsp_xbar_demux_002_src2_valid;                                                                     // rsp_xbar_demux_002:src2_valid -> width_adapter_011:in_valid
	wire          rsp_xbar_demux_002_src2_startofpacket;                                                             // rsp_xbar_demux_002:src2_startofpacket -> width_adapter_011:in_startofpacket
	wire   [88:0] rsp_xbar_demux_002_src2_data;                                                                      // rsp_xbar_demux_002:src2_data -> width_adapter_011:in_data
	wire   [15:0] rsp_xbar_demux_002_src2_channel;                                                                   // rsp_xbar_demux_002:src2_channel -> width_adapter_011:in_channel
	wire          rsp_xbar_demux_002_src2_ready;                                                                     // width_adapter_011:in_ready -> rsp_xbar_demux_002:src2_ready
	wire          width_adapter_011_src_endofpacket;                                                                 // width_adapter_011:out_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          width_adapter_011_src_valid;                                                                       // width_adapter_011:out_valid -> rsp_xbar_mux_002:sink1_valid
	wire          width_adapter_011_src_startofpacket;                                                               // width_adapter_011:out_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [106:0] width_adapter_011_src_data;                                                                        // width_adapter_011:out_data -> rsp_xbar_mux_002:sink1_data
	wire          width_adapter_011_src_ready;                                                                       // rsp_xbar_mux_002:sink1_ready -> width_adapter_011:out_ready
	wire   [15:0] width_adapter_011_src_channel;                                                                     // width_adapter_011:out_channel -> rsp_xbar_mux_002:sink1_channel
	wire          crosser_out_endofpacket;                                                                           // crosser:out_endofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_out_valid;                                                                                 // crosser:out_valid -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_out_startofpacket;                                                                         // crosser:out_startofpacket -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] crosser_out_data;                                                                                  // crosser:out_data -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [15:0] crosser_out_channel;                                                                               // crosser:out_channel -> altpll_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                               // cmd_xbar_demux_001:src6_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                     // cmd_xbar_demux_001:src6_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                             // cmd_xbar_demux_001:src6_startofpacket -> crosser:in_startofpacket
	wire  [106:0] cmd_xbar_demux_001_src6_data;                                                                      // cmd_xbar_demux_001:src6_data -> crosser:in_data
	wire   [15:0] cmd_xbar_demux_001_src6_channel;                                                                   // cmd_xbar_demux_001:src6_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src6_ready;                                                                     // crosser:in_ready -> cmd_xbar_demux_001:src6_ready
	wire          crosser_001_out_endofpacket;                                                                       // crosser_001:out_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          crosser_001_out_valid;                                                                             // crosser_001:out_valid -> rsp_xbar_mux_001:sink6_valid
	wire          crosser_001_out_startofpacket;                                                                     // crosser_001:out_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [106:0] crosser_001_out_data;                                                                              // crosser_001:out_data -> rsp_xbar_mux_001:sink6_data
	wire   [15:0] crosser_001_out_channel;                                                                           // crosser_001:out_channel -> rsp_xbar_mux_001:sink6_channel
	wire          crosser_001_out_ready;                                                                             // rsp_xbar_mux_001:sink6_ready -> crosser_001:out_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                               // rsp_xbar_demux_006:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                     // rsp_xbar_demux_006:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                             // rsp_xbar_demux_006:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [106:0] rsp_xbar_demux_006_src0_data;                                                                      // rsp_xbar_demux_006:src0_data -> crosser_001:in_data
	wire   [15:0] rsp_xbar_demux_006_src0_channel;                                                                   // rsp_xbar_demux_006:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                     // crosser_001:in_ready -> rsp_xbar_demux_006:src0_ready
	wire   [15:0] limiter_cmd_valid_data;                                                                            // limiter:cmd_src_valid -> cmd_xbar_demux_002:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                          // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                          // epcs_flash:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                          // systimer:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                          // timestamp:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                          // uart1:irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                                                          // uart2:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                                                          // uart3:irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver7_irq;                                                                          // pio_key:irq -> irq_mapper:receiver7_irq
	wire          irq_mapper_receiver8_irq;                                                                          // oc_i2c_master_0:wb_inta_o -> irq_mapper:receiver8_irq
	wire          irq_mapper_receiver9_irq;                                                                          // dma_0:dma_ctl_irq -> irq_mapper:receiver9_irq
	wire   [31:0] nios2_d_irq_irq;                                                                                   // irq_mapper:sender_irq -> nios2:d_irq

	nios2_nios2 nios2 (
		.clk                                   (altpll_c0_clk),                                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                    //                   reset_n.reset_n
		.d_address                             (nios2_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_data_master_writedata),                                        //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                               //                          .waitrequest
		.d_irq                                 (nios2_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                    // custom_instruction_master.readra
	);

	nios2_onchip_ram onchip_ram (
		.clk        (altpll_c0_clk),                                           //   clk1.clk
		.address    (onchip_ram_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_ram_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_ram_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_ram_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_ram_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_ram_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_ram_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                           // reset1.reset
	);

	nios2_sysid sysid (
		.clock    (altpll_c0_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                             //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	nios2_jtag_uart jtag_uart (
		.clk            (altpll_c0_clk),                                                          //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	nios2_sdram sdram (
		.clk            (altpll_c0_clk),                                         //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                       // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                            //  wire.export
		.zs_ba          (sdram_ba),                                              //      .export
		.zs_cas_n       (sdram_cas_n),                                           //      .export
		.zs_cke         (sdram_cke),                                             //      .export
		.zs_cs_n        (sdram_cs_n),                                            //      .export
		.zs_dq          (sdram_dq),                                              //      .export
		.zs_dqm         (sdram_dqm),                                             //      .export
		.zs_ras_n       (sdram_ras_n),                                           //      .export
		.zs_we_n        (sdram_we_n)                                             //      .export
	);

	nios2_epcs_flash epcs_flash (
		.clk           (altpll_c0_clk),                                                          //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.address       (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_address),    // epcs_control_port.address
		.chipselect    (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_chipselect), //                  .chipselect
		.dataavailable (),                                                                       //                  .dataavailable
		.endofpacket   (),                                                                       //                  .endofpacket
		.read_n        (~epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_read),      //                  .read_n
		.readdata      (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_readdata),   //                  .readdata
		.readyfordata  (),                                                                       //                  .readyfordata
		.write_n       (~epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_write),     //                  .write_n
		.writedata     (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver1_irq)                                                //               irq.irq
	);

	nios2_altpll altpll (
		.clk       (clk_clk),                                                   //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),                        // inclk_interface_reset.reset
		.read      (altpll_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (altpll_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (altpll_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (altpll_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (altpll_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (altpll_c0_clk),                                             //                    c0.clk
		.c1        (sdram_clk_clk),                                             //                    c1.clk
		.areset    (),                                                          //        areset_conduit.export
		.locked    (),                                                          //        locked_conduit.export
		.phasedone ()                                                           //     phasedone_conduit.export
	);

	nios2_systimer systimer (
		.clk        (altpll_c0_clk),                                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       // reset.reset_n
		.address    (systimer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (systimer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (systimer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (systimer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~systimer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                               //   irq.irq
	);

	nios2_timestamp timestamp (
		.clk        (altpll_c0_clk),                                          //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        // reset.reset_n
		.address    (timestamp_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timestamp_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timestamp_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timestamp_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timestamp_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                                //   irq.irq
	);

	nios2_uart1 uart1 (
		.clk           (altpll_c0_clk),                                         //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address       (uart1_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart1_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart1_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart1_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart1_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart1_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart1_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                      //                    .dataavailable
		.readyfordata  (),                                                      //                    .readyfordata
		.rxd           (uart1_rxd),                                             // external_connection.export
		.txd           (uart1_txd),                                             //                    .export
		.irq           (irq_mapper_receiver4_irq)                               //                 irq.irq
	);

	nios2_uart1 uart2 (
		.clk           (altpll_c0_clk),                                         //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address       (uart2_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart2_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart2_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart2_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart2_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart2_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart2_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                      //                    .dataavailable
		.readyfordata  (),                                                      //                    .readyfordata
		.rxd           (uart2_rxd),                                             // external_connection.export
		.txd           (uart2_txd),                                             //                    .export
		.irq           (irq_mapper_receiver5_irq)                               //                 irq.irq
	);

	nios2_uart1 uart3 (
		.clk           (altpll_c0_clk),                                         //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address       (uart3_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart3_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart3_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart3_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart3_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart3_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart3_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                      //                    .dataavailable
		.readyfordata  (),                                                      //                    .readyfordata
		.rxd           (uart3_rxd),                                             // external_connection.export
		.txd           (uart3_txd),                                             //                    .export
		.irq           (irq_mapper_receiver6_irq)                               //                 irq.irq
	);

	nios2_pio_led pio_led (
		.clk        (altpll_c0_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (pio_led_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_led_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_led_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_led_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_led_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_export)                                            // external_connection.export
	);

	nios2_pio_key pio_key (
		.clk        (altpll_c0_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (pio_key_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_key_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_key_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_key_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_key_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (key_export),                                           // external_connection.export
		.irq        (irq_mapper_receiver7_irq)                              //                 irq.irq
	);

	oc_i2c_master oc_i2c_master_0 (
		.wb_clk_i   (altpll_c0_clk),                                                   //       s1_clk.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                  // s1_clk_reset.reset
		.wb_ack_o   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_waitrequest),   //           s1.waitrequest_n
		.wb_adr_i   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_address),       //             .address
		.wb_dat_i   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_writedata),     //             .writedata
		.wb_dat_o   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_readdata),      //             .readdata
		.wb_stb_i   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_begintransfer), //             .begintransfer
		.wb_we_i    (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_write),         //             .write
		.wb_cyc_i   (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_chipselect),    //             .chipselect
		.scl_pad_io (oc_i2c_master_scl_pad_io),                                        //       global.export
		.sda_pad_io (oc_i2c_master_sda_pad_io),                                        //             .export
		.wb_inta_o  (irq_mapper_receiver8_irq)                                         //       s1_irq.irq
	);

	nios2_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (altpll_c0_clk),                      //          clk.clk
		.clk_reset_reset      (rst_controller_002_reset_out_reset), //    clk_reset.reset
		.master_address       (master_0_master_address),            //       master.address
		.master_readdata      (master_0_master_readdata),           //             .readdata
		.master_read          (master_0_master_read),               //             .read
		.master_write         (master_0_master_write),              //             .write
		.master_writedata     (master_0_master_writedata),          //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),        //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid),      //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),         //             .byteenable
		.master_reset_reset   ()                                    // master_reset.reset
	);

	nios2_dma_0 dma_0 (
		.clk                (altpll_c0_clk),                                                      //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                                    //              reset.reset_n
		.dma_ctl_address    (dma_0_control_port_slave_translator_avalon_anti_slave_0_address),    // control_port_slave.address
		.dma_ctl_chipselect (dma_0_control_port_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.dma_ctl_readdata   (dma_0_control_port_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.dma_ctl_write_n    (~dma_0_control_port_slave_translator_avalon_anti_slave_0_write),     //                   .write_n
		.dma_ctl_writedata  (dma_0_control_port_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver9_irq),                                           //                irq.irq
		.read_address       (dma_0_read_master_address),                                          //        read_master.address
		.read_chipselect    (dma_0_read_master_chipselect),                                       //                   .chipselect
		.read_read_n        (dma_0_read_master_read),                                             //                   .read_n
		.read_readdata      (dma_0_read_master_readdata),                                         //                   .readdata
		.read_readdatavalid (dma_0_read_master_readdatavalid),                                    //                   .readdatavalid
		.read_waitrequest   (dma_0_read_master_waitrequest),                                      //                   .waitrequest
		.write_address      (dma_0_write_master_address),                                         //       write_master.address
		.write_chipselect   (dma_0_write_master_chipselect),                                      //                   .chipselect
		.write_waitrequest  (dma_0_write_master_waitrequest),                                     //                   .waitrequest
		.write_write_n      (dma_0_write_master_write),                                           //                   .write_n
		.write_writedata    (dma_0_write_master_writedata),                                       //                   .writedata
		.write_byteenable   (dma_0_write_master_byteenable)                                       //                   .byteenable
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_instruction_master_translator (
		.clk                      (altpll_c0_clk),                                                               //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_instruction_master_readdata),                                           //                          .readdata
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_byteenable            (4'b1111),                                                                     //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                            //               (terminated)
		.av_write                 (1'b0),                                                                        //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.av_debugaccess           (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (1)
	) nios2_data_master_translator (
		.clk                      (altpll_c0_clk),                                                        //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address              (nios2_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_data_master_read),                                               //                          .read
		.av_readdata              (nios2_data_master_readdata),                                           //                          .readdata
		.av_write                 (nios2_data_master_write),                                              //                          .write
		.av_writedata             (nios2_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                 //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_chipselect            (1'b0),                                                                 //               (terminated)
		.av_readdatavalid         (),                                                                     //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) master_0_master_translator (
		.clk                      (altpll_c0_clk),                                                      //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                     //                     reset.reset
		.uav_address              (master_0_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (master_0_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (master_0_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (master_0_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (master_0_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (master_0_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (master_0_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (master_0_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (master_0_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (master_0_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (master_0_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (master_0_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (master_0_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (master_0_master_byteenable),                                         //                          .byteenable
		.av_read                  (master_0_master_read),                                               //                          .read
		.av_readdata              (master_0_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (master_0_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (master_0_master_write),                                              //                          .write
		.av_writedata             (master_0_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                               //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (25),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_0_write_master_translator (
		.clk                      (altpll_c0_clk),                                                         //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                     reset.reset
		.uav_address              (dma_0_write_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_0_write_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_0_write_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_0_write_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_0_write_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_0_write_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_0_write_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_0_write_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_0_write_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_0_write_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_0_write_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_0_write_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_0_write_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (dma_0_write_master_byteenable),                                         //                          .byteenable
		.av_chipselect            (dma_0_write_master_chipselect),                                         //                          .chipselect
		.av_write                 (~dma_0_write_master_write),                                             //                          .write
		.av_writedata             (dma_0_write_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                  //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                  //               (terminated)
		.av_begintransfer         (1'b0),                                                                  //               (terminated)
		.av_read                  (1'b0),                                                                  //               (terminated)
		.av_readdata              (),                                                                      //               (terminated)
		.av_readdatavalid         (),                                                                      //               (terminated)
		.av_lock                  (1'b0),                                                                  //               (terminated)
		.av_debugaccess           (1'b0),                                                                  //               (terminated)
		.uav_clken                (),                                                                      //               (terminated)
		.av_clken                 (1'b1),                                                                  //               (terminated)
		.uav_response             (2'b00),                                                                 //               (terminated)
		.av_response              (),                                                                      //               (terminated)
		.uav_writeresponserequest (),                                                                      //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                  //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                  //               (terminated)
		.av_writeresponsevalid    ()                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (24),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_0_read_master_translator (
		.clk                      (altpll_c0_clk),                                                        //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                       //                     reset.reset
		.uav_address              (dma_0_read_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_0_read_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_0_read_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_0_read_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_0_read_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_0_read_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_0_read_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_0_read_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_0_read_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_0_read_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_0_read_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_0_read_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_0_read_master_waitrequest),                                        //                          .waitrequest
		.av_chipselect            (dma_0_read_master_chipselect),                                         //                          .chipselect
		.av_read                  (~dma_0_read_master_read),                                              //                          .read
		.av_readdata              (dma_0_read_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (dma_0_read_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                 //               (terminated)
		.av_byteenable            (2'b11),                                                                //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                 //               (terminated)
		.av_begintransfer         (1'b0),                                                                 //               (terminated)
		.av_write                 (1'b0),                                                                 //               (terminated)
		.av_writedata             (16'b0000000000000000),                                                 //               (terminated)
		.av_lock                  (1'b0),                                                                 //               (terminated)
		.av_debugaccess           (1'b0),                                                                 //               (terminated)
		.uav_clken                (),                                                                     //               (terminated)
		.av_clken                 (1'b1),                                                                 //               (terminated)
		.uav_response             (2'b00),                                                                //               (terminated)
		.av_response              (),                                                                     //               (terminated)
		.uav_writeresponserequest (),                                                                     //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                 //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                 //               (terminated)
		.av_writeresponsevalid    ()                                                                      //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_jtag_debug_module_translator (
		.clk                      (altpll_c0_clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_chipselect            (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (11),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_ram_s1_translator (
		.clk                      (altpll_c0_clk),                                                            //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address              (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_ram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_ram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_ram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_ram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_ram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_ram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_ram_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (altpll_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) epcs_flash_epcs_control_port_translator (
		.clk                      (altpll_c0_clk),                                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address              (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (epcs_flash_epcs_control_port_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                                        //              (terminated)
		.av_burstcount            (),                                                                                        //              (terminated)
		.av_byteenable            (),                                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                        //              (terminated)
		.av_lock                  (),                                                                                        //              (terminated)
		.av_clken                 (),                                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                                    //              (terminated)
		.av_debugaccess           (),                                                                                        //              (terminated)
		.av_outputenable          (),                                                                                        //              (terminated)
		.uav_response             (),                                                                                        //              (terminated)
		.av_response              (2'b00),                                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (altpll_c0_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (altpll_c0_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altpll_pll_slave_translator (
		.clk                      (clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                          //                    reset.reset
		.uav_address              (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (altpll_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (altpll_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (altpll_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (altpll_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (altpll_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_chipselect            (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) systimer_s1_translator (
		.clk                      (altpll_c0_clk),                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address              (systimer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (systimer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (systimer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (systimer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (systimer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (systimer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (systimer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (systimer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (systimer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (systimer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (systimer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (systimer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (systimer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (systimer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                       //              (terminated)
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                       //              (terminated)
		.av_burstcount            (),                                                                       //              (terminated)
		.av_byteenable            (),                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                   //              (terminated)
		.av_waitrequest           (1'b0),                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timestamp_s1_translator (
		.clk                      (altpll_c0_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address              (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timestamp_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timestamp_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timestamp_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timestamp_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timestamp_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart1_s1_translator (
		.clk                      (altpll_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (uart1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (uart1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (uart1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (uart1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (uart1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (uart1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (uart1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (uart1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (uart1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (uart1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (uart1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (uart1_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (uart1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (uart1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (uart1_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (uart1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart2_s1_translator (
		.clk                      (altpll_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (uart2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (uart2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (uart2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (uart2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (uart2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (uart2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (uart2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (uart2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (uart2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (uart2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (uart2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (uart2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (uart2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (uart2_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (uart2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (uart2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (uart2_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (uart2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart3_s1_translator (
		.clk                      (altpll_c0_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (uart3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (uart3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (uart3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (uart3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (uart3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (uart3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (uart3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (uart3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (uart3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (uart3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (uart3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (uart3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (uart3_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (uart3_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (uart3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (uart3_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (uart3_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect            (uart3_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_led_s1_translator (
		.clk                      (altpll_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_led_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_led_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_led_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_led_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_led_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_key_s1_translator (
		.clk                      (altpll_c0_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_key_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_key_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_key_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_key_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_key_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) oc_i2c_master_0_s1_translator (
		.clk                      (altpll_c0_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address              (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_waitrequest           (~oc_i2c_master_0_s1_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_chipselect            (oc_i2c_master_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                              //              (terminated)
		.av_beginbursttransfer    (),                                                                              //              (terminated)
		.av_burstcount            (),                                                                              //              (terminated)
		.av_byteenable            (),                                                                              //              (terminated)
		.av_readdatavalid         (1'b0),                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                              //              (terminated)
		.av_lock                  (),                                                                              //              (terminated)
		.av_clken                 (),                                                                              //              (terminated)
		.uav_clken                (1'b0),                                                                          //              (terminated)
		.av_debugaccess           (),                                                                              //              (terminated)
		.av_outputenable          (),                                                                              //              (terminated)
		.uav_response             (),                                                                              //              (terminated)
		.av_response              (2'b00),                                                                         //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                          //              (terminated)
		.uav_writeresponsevalid   (),                                                                              //              (terminated)
		.av_writeresponserequest  (),                                                                              //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dma_0_control_port_slave_translator (
		.clk                      (altpll_c0_clk),                                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address              (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dma_0_control_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dma_0_control_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (dma_0_control_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dma_0_control_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (dma_0_control_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                    //              (terminated)
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_byteenable            (),                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (4),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (altpll_c0_clk),                                                                        //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_src_valid),                                                               //        rp.valid
		.rp_data                 (rsp_xbar_mux_src_data),                                                                //          .data
		.rp_channel              (rsp_xbar_mux_src_channel),                                                             //          .channel
		.rp_startofpacket        (rsp_xbar_mux_src_startofpacket),                                                       //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_src_endofpacket),                                                         //          .endofpacket
		.rp_ready                (rsp_xbar_mux_src_ready),                                                               //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (altpll_c0_clk),                                                                 //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address              (nios2_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_001_src_valid),                                                    //        rp.valid
		.rp_data                 (rsp_xbar_mux_001_src_data),                                                     //          .data
		.rp_channel              (rsp_xbar_mux_001_src_channel),                                                  //          .channel
		.rp_startofpacket        (rsp_xbar_mux_001_src_startofpacket),                                            //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_001_src_endofpacket),                                              //          .endofpacket
		.rp_ready                (rsp_xbar_mux_001_src_ready),                                                    //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) master_0_master_translator_avalon_universal_master_0_agent (
		.clk                     (altpll_c0_clk),                                                               //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.av_address              (master_0_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (master_0_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (master_0_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (master_0_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (master_0_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (master_0_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (master_0_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (master_0_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (master_0_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (master_0_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (master_0_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (master_0_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (master_0_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (master_0_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                       //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                        //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                     //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                 //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                       //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (75),
		.PKT_THREAD_ID_H           (79),
		.PKT_THREAD_ID_L           (79),
		.PKT_CACHE_H               (86),
		.PKT_CACHE_L               (83),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_0_read_master_translator_avalon_universal_master_0_agent (
		.clk                     (altpll_c0_clk),                                                                 //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.av_address              (dma_0_read_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_0_read_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_0_read_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_0_read_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_0_read_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_0_read_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_0_read_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_0_read_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_0_read_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_0_read_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_0_read_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_002_src3_valid),                                                 //        rp.valid
		.rp_data                 (rsp_xbar_demux_002_src3_data),                                                  //          .data
		.rp_channel              (rsp_xbar_demux_002_src3_channel),                                               //          .channel
		.rp_startofpacket        (rsp_xbar_demux_002_src3_startofpacket),                                         //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_002_src3_endofpacket),                                           //          .endofpacket
		.rp_ready                (rsp_xbar_demux_002_src3_ready),                                                 //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (75),
		.PKT_THREAD_ID_H           (79),
		.PKT_THREAD_ID_L           (79),
		.PKT_CACHE_H               (86),
		.PKT_CACHE_L               (83),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (16),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_0_write_master_translator_avalon_universal_master_0_agent (
		.clk                     (altpll_c0_clk),                                                                  //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.av_address              (dma_0_write_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_0_write_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_0_write_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_0_write_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_0_write_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_0_write_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_0_write_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_0_write_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_0_write_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_0_write_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_0_write_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_001_src3_valid),                                                  //        rp.valid
		.rp_data                 (rsp_xbar_demux_001_src3_data),                                                   //          .data
		.rp_channel              (rsp_xbar_demux_001_src3_channel),                                                //          .channel
		.rp_startofpacket        (rsp_xbar_demux_001_src3_startofpacket),                                          //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_001_src3_endofpacket),                                            //          .endofpacket
		.rp_ready                (rsp_xbar_demux_001_src3_ready),                                                  //          .ready
		.av_response             (),                                                                               // (terminated)
		.av_writeresponserequest (1'b0),                                                                           // (terminated)
		.av_writeresponsevalid   ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                       //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                       //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                        //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                     //                .channel
		.rf_sink_ready           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_ram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                      //                .channel
		.rf_sink_ready           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (74),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (78),
		.PKT_DEST_ID_L             (75),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (82),
		.PKT_PROTECTION_L          (80),
		.PKT_RESPONSE_STATUS_H     (88),
		.PKT_RESPONSE_STATUS_L     (87),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (89),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                               //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                               //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                         //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                             //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (90),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (altpll_c0_clk),                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                                        //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                                        //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                                         //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                                      //                .channel
		.rf_sink_ready           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) altpll_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altpll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_out_ready),                                                                     //              cp.ready
		.cp_valid                (crosser_out_valid),                                                                     //                .valid
		.cp_data                 (crosser_out_data),                                                                      //                .data
		.cp_startofpacket        (crosser_out_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (crosser_out_endofpacket),                                                               //                .endofpacket
		.cp_channel              (crosser_out_channel),                                                                   //                .channel
		.rf_sink_ready           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                              // clk_reset.reset
		.in_data           (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_startofpacket  (1'b0),                                                                            // (terminated)
		.in_endofpacket    (1'b0),                                                                            // (terminated)
		.out_startofpacket (),                                                                                // (terminated)
		.out_endofpacket   (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) systimer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (systimer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (systimer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (systimer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (systimer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (systimer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (systimer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (systimer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (systimer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (systimer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (systimer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (systimer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (systimer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (systimer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (systimer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (systimer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                  //                .channel
		.rf_sink_ready           (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (systimer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (systimer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (systimer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timestamp_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timestamp_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                   //                .channel
		.rf_sink_ready           (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timestamp_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timestamp_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) uart1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (uart1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                               //                .channel
		.rf_sink_ready           (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) uart2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (uart2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_010_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_010_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_010_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_010_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_010_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_010_src_channel),                                                  //                .channel
		.rf_sink_ready           (uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) uart3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (uart3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                              //                .channel
		.rf_sink_ready           (uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_led_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_led_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                //                .channel
		.rf_sink_ready           (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_led_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_led_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_key_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_key_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                //                .channel
		.rf_sink_ready           (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_key_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_key_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_key_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src14_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src14_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src14_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src14_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src14_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src14_channel),                                                        //                .channel
		.rf_sink_ready           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                   //     (terminated)
		.m0_writeresponserequest (),                                                                                        //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                     //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (16),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_0_control_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (altpll_c0_clk),                                                                                 //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_015_src_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_015_src_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_015_src_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_015_src_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_015_src_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_015_src_channel),                                                                  //                .channel
		.rf_sink_ready           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (altpll_c0_clk),                                                                                 //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	nios2_addr_router addr_router (
		.sink_ready         (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                //       src.ready
		.src_valid          (addr_router_src_valid),                                                                //          .valid
		.src_data           (addr_router_src_data),                                                                 //          .data
		.src_channel        (addr_router_src_channel),                                                              //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                           //          .endofpacket
	);

	nios2_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                     //          .valid
		.src_data           (addr_router_001_src_data),                                                      //          .data
		.src_channel        (addr_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                //          .endofpacket
	);

	nios2_addr_router_002 addr_router_002 (
		.sink_ready         (master_0_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (master_0_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (master_0_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                   //          .valid
		.src_data           (addr_router_002_src_data),                                                    //          .data
		.src_channel        (addr_router_002_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                              //          .endofpacket
	);

	nios2_addr_router_003 addr_router_003 (
		.sink_ready         (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                     //          .valid
		.src_data           (addr_router_003_src_data),                                                      //          .data
		.src_channel        (addr_router_003_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                                //          .endofpacket
	);

	nios2_addr_router_004 addr_router_004 (
		.sink_ready         (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                      //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                      //          .valid
		.src_data           (addr_router_004_src_data),                                                       //          .data
		.src_channel        (addr_router_004_src_channel),                                                    //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                 //          .endofpacket
	);

	nios2_id_router id_router (
		.sink_ready         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                //       src.ready
		.src_valid          (id_router_src_valid),                                                                //          .valid
		.src_data           (id_router_src_data),                                                                 //          .data
		.src_channel        (id_router_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                           //          .endofpacket
	);

	nios2_id_router_001 id_router_001 (
		.sink_ready         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_ram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                  //       src.ready
		.src_valid          (id_router_001_src_valid),                                                  //          .valid
		.src_data           (id_router_001_src_data),                                                   //          .data
		.src_channel        (id_router_001_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                             //          .endofpacket
	);

	nios2_id_router_002 id_router_002 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                             //       src.ready
		.src_valid          (id_router_002_src_valid),                                             //          .valid
		.src_data           (id_router_002_src_data),                                              //          .data
		.src_channel        (id_router_002_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                        //          .endofpacket
	);

	nios2_id_router id_router_003 (
		.sink_ready         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (epcs_flash_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                 //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                 //          .valid
		.src_data           (id_router_003_src_data),                                                                  //          .data
		.src_channel        (id_router_003_src_channel),                                                               //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                         //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                            //          .endofpacket
	);

	nios2_id_router_004 id_router_004 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                        //       src.ready
		.src_valid          (id_router_004_src_valid),                                                        //          .valid
		.src_data           (id_router_004_src_data),                                                         //          .data
		.src_channel        (id_router_004_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                   //          .endofpacket
	);

	nios2_id_router_004 id_router_005 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                //          .valid
		.src_data           (id_router_005_src_data),                                                                 //          .data
		.src_channel        (id_router_005_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                           //          .endofpacket
	);

	nios2_id_router_004 id_router_006 (
		.sink_ready         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altpll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                     //       src.ready
		.src_valid          (id_router_006_src_valid),                                                     //          .valid
		.src_data           (id_router_006_src_data),                                                      //          .data
		.src_channel        (id_router_006_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                //          .endofpacket
	);

	nios2_id_router_004 id_router_007 (
		.sink_ready         (systimer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (systimer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (systimer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (systimer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (systimer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                //       src.ready
		.src_valid          (id_router_007_src_valid),                                                //          .valid
		.src_data           (id_router_007_src_data),                                                 //          .data
		.src_channel        (id_router_007_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                           //          .endofpacket
	);

	nios2_id_router_004 id_router_008 (
		.sink_ready         (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timestamp_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                 //       src.ready
		.src_valid          (id_router_008_src_valid),                                                 //          .valid
		.src_data           (id_router_008_src_data),                                                  //          .data
		.src_channel        (id_router_008_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                            //          .endofpacket
	);

	nios2_id_router_004 id_router_009 (
		.sink_ready         (uart1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                             //       src.ready
		.src_valid          (id_router_009_src_valid),                                             //          .valid
		.src_data           (id_router_009_src_data),                                              //          .data
		.src_channel        (id_router_009_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                        //          .endofpacket
	);

	nios2_id_router_010 id_router_010 (
		.sink_ready         (uart2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                             //       src.ready
		.src_valid          (id_router_010_src_valid),                                             //          .valid
		.src_data           (id_router_010_src_data),                                              //          .data
		.src_channel        (id_router_010_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                        //          .endofpacket
	);

	nios2_id_router_004 id_router_011 (
		.sink_ready         (uart3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                             //       src.ready
		.src_valid          (id_router_011_src_valid),                                             //          .valid
		.src_data           (id_router_011_src_data),                                              //          .data
		.src_channel        (id_router_011_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                        //          .endofpacket
	);

	nios2_id_router_004 id_router_012 (
		.sink_ready         (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_led_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                               //       src.ready
		.src_valid          (id_router_012_src_valid),                                               //          .valid
		.src_data           (id_router_012_src_data),                                                //          .data
		.src_channel        (id_router_012_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                          //          .endofpacket
	);

	nios2_id_router_004 id_router_013 (
		.sink_ready         (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_key_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                               //       src.ready
		.src_valid          (id_router_013_src_valid),                                               //          .valid
		.src_data           (id_router_013_src_data),                                                //          .data
		.src_channel        (id_router_013_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                          //          .endofpacket
	);

	nios2_id_router_004 id_router_014 (
		.sink_ready         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (oc_i2c_master_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                       //       src.ready
		.src_valid          (id_router_014_src_valid),                                                       //          .valid
		.src_data           (id_router_014_src_data),                                                        //          .data
		.src_channel        (id_router_014_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                  //          .endofpacket
	);

	nios2_id_router_010 id_router_015 (
		.sink_ready         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (altpll_c0_clk),                                                                       //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                             //       src.ready
		.src_valid          (id_router_015_src_valid),                                                             //          .valid
		.src_data           (id_router_015_src_data),                                                              //          .data
		.src_channel        (id_router_015_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                        //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (93),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (16),
		.VALID_WIDTH               (16),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (altpll_c0_clk),                      //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_002_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_002_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_002_src_data),           //          .data
		.cmd_sink_channel       (addr_router_002_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_002_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_002_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_002_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_002_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_002_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_002_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_002_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (16),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (altpll_c0_clk),                       //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_001_src_valid),          //     sink0.valid
		.sink0_data            (cmd_xbar_mux_001_src_data),           //          .data
		.sink0_channel         (cmd_xbar_mux_001_src_channel),        //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_001_src_startofpacket),  //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_001_src_endofpacket),    //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_001_src_ready),          //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (89),
		.ST_CHANNEL_W              (16),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (altpll_c0_clk),                           //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_002_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_002_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_002_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_002_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_002_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_002_src_ready),              //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (altpll_c0_clk),                       //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                      // reset_in0.reset
		.reset_in1  (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                             //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("none"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (nios2_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1  (~reset_reset_n),                      // reset_in1.reset
		.clk        (),                                    //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset),  // reset_out.reset
		.reset_in2  (1'b0),                                // (terminated)
		.reset_in3  (1'b0),                                // (terminated)
		.reset_in4  (1'b0),                                // (terminated)
		.reset_in5  (1'b0),                                // (terminated)
		.reset_in6  (1'b0),                                // (terminated)
		.reset_in7  (1'b0),                                // (terminated)
		.reset_in8  (1'b0),                                // (terminated)
		.reset_in9  (1'b0),                                // (terminated)
		.reset_in10 (1'b0),                                // (terminated)
		.reset_in11 (1'b0),                                // (terminated)
		.reset_in12 (1'b0),                                // (terminated)
		.reset_in13 (1'b0),                                // (terminated)
		.reset_in14 (1'b0),                                // (terminated)
		.reset_in15 (1'b0)                                 // (terminated)
	);

	nios2_cmd_xbar_demux cmd_xbar_demux (
		.clk                (altpll_c0_clk),                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_src_ready),             //      sink.ready
		.sink_channel       (addr_router_src_channel),           //          .channel
		.sink_data          (addr_router_src_data),              //          .data
		.sink_startofpacket (addr_router_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //      src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //          .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //          .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //          .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //          .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //      src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //          .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //          .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //          .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (altpll_c0_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.sink_ready          (addr_router_001_src_ready),              //      sink.ready
		.sink_channel        (addr_router_001_src_channel),            //          .channel
		.sink_data           (addr_router_001_src_data),               //          .data
		.sink_startofpacket  (addr_router_001_src_startofpacket),      //          .startofpacket
		.sink_endofpacket    (addr_router_001_src_endofpacket),        //          .endofpacket
		.sink_valid          (addr_router_001_src_valid),              //          .valid
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //      src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //          .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //          .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //          .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //          .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //      src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //          .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //          .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //          .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //          .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //          .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //      src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //          .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //          .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //          .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //          .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //          .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //      src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //          .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //          .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //          .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //          .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //          .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //      src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //          .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //          .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //          .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //          .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //          .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //      src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //          .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //          .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //          .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //          .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //          .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //      src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //          .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //          .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //          .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //          .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //          .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //      src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //          .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //          .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //          .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //          .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //          .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //      src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //          .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //          .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //          .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //          .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //          .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //      src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //          .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //          .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //          .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //          .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //          .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //     src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //     src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //          .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //     src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //          .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //     src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //          .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //     src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //          .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //     src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (altpll_c0_clk),                         //        clk.clk
		.reset              (rst_controller_reset_out_reset),        //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),                 //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),               //           .channel
		.sink_data          (limiter_cmd_src_data),                  //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),         //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),           //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),                // sink_valid.data
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_002_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_002_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_002_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_002_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_002_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_002_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_002_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_002_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_002_src3_endofpacket)    //           .endofpacket
	);

	nios2_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_demux_003 cmd_xbar_demux_004 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (altpll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (altpll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_src_ready),               //     sink0.ready
		.sink0_valid         (width_adapter_src_valid),               //          .valid
		.sink0_channel       (width_adapter_src_channel),             //          .channel
		.sink0_data          (width_adapter_src_data),                //          .data
		.sink0_startofpacket (width_adapter_src_startofpacket),       //          .startofpacket
		.sink0_endofpacket   (width_adapter_src_endofpacket),         //          .endofpacket
		.sink1_ready         (width_adapter_002_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_002_src_valid),           //          .valid
		.sink1_channel       (width_adapter_002_src_channel),         //          .channel
		.sink1_data          (width_adapter_002_src_data),            //          .data
		.sink1_startofpacket (width_adapter_002_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_002_src_endofpacket),     //          .endofpacket
		.sink2_ready         (width_adapter_004_src_ready),           //     sink2.ready
		.sink2_valid         (width_adapter_004_src_valid),           //          .valid
		.sink2_channel       (width_adapter_004_src_channel),         //          .channel
		.sink2_data          (width_adapter_004_src_data),            //          .data
		.sink2_startofpacket (width_adapter_004_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket   (width_adapter_004_src_endofpacket),     //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_004_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_mux_001 cmd_xbar_mux_002 (
		.clk                 (altpll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_001_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_001_src_valid),           //          .valid
		.sink0_channel       (width_adapter_001_src_channel),         //          .channel
		.sink0_data          (width_adapter_001_src_data),            //          .data
		.sink0_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink1_ready         (width_adapter_003_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_003_src_valid),           //          .valid
		.sink1_channel       (width_adapter_003_src_channel),         //          .channel
		.sink1_data          (width_adapter_003_src_data),            //          .data
		.sink1_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink2_ready         (width_adapter_005_src_ready),           //     sink2.ready
		.sink2_valid         (width_adapter_005_src_valid),           //          .valid
		.sink2_channel       (width_adapter_005_src_channel),         //          .channel
		.sink2_data          (width_adapter_005_src_data),            //          .data
		.sink2_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink3_ready         (cmd_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_mux cmd_xbar_mux_003 (
		.clk                 (altpll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src3_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src3_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src3_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src3_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src3_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src3_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	nios2_cmd_xbar_mux cmd_xbar_mux_010 (
		.clk                 (altpll_c0_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src10_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src2_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src2_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src2_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_002_src2_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src2_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src2_endofpacket)     //          .endofpacket
	);

	nios2_cmd_xbar_mux cmd_xbar_mux_015 (
		.clk                 (altpll_c0_clk),                          //       clk.clk
		.reset               (rst_controller_reset_out_reset),         // clk_reset.reset
		.src_ready           (cmd_xbar_mux_015_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_015_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_015_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_015_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_015_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_015_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src15_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src15_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src15_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src15_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src3_ready),          //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src3_valid),          //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src3_channel),        //          .channel
		.sink1_data          (cmd_xbar_demux_002_src3_data),           //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src3_startofpacket),  //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src3_endofpacket)     //          .endofpacket
	);

	nios2_rsp_xbar_demux rsp_xbar_demux (
		.clk                (altpll_c0_clk),                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_001_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_001_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_001_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_001_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_001_src3_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_001 rsp_xbar_demux_002 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_002_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_002_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_002_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_002_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.src3_ready         (rsp_xbar_demux_002_src3_ready),         //      src3.ready
		.src3_valid         (rsp_xbar_demux_002_src3_valid),         //          .valid
		.src3_data          (rsp_xbar_demux_002_src3_data),          //          .data
		.src3_channel       (rsp_xbar_demux_002_src3_channel),       //          .channel
		.src3_startofpacket (rsp_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.src3_endofpacket   (rsp_xbar_demux_002_src3_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_004 rsp_xbar_demux_004 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_004 rsp_xbar_demux_005 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_004 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_004 rsp_xbar_demux_007 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_004 rsp_xbar_demux_008 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_004 rsp_xbar_demux_009 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux rsp_xbar_demux_010 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_004 rsp_xbar_demux_011 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_004 rsp_xbar_demux_012 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_004 rsp_xbar_demux_013 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux_004 rsp_xbar_demux_014 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_demux rsp_xbar_demux_015 (
		.clk                (altpll_c0_clk),                         //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_015_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_015_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_015_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_015_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_015_src1_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (altpll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (width_adapter_006_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_006_src_valid),           //          .valid
		.sink1_channel       (width_adapter_006_src_channel),         //          .channel
		.sink1_data          (width_adapter_006_src_data),            //          .data
		.sink1_startofpacket (width_adapter_006_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_006_src_endofpacket),     //          .endofpacket
		.sink2_ready         (width_adapter_009_src_ready),           //     sink2.ready
		.sink2_valid         (width_adapter_009_src_valid),           //          .valid
		.sink2_channel       (width_adapter_009_src_channel),         //          .channel
		.sink2_data          (width_adapter_009_src_data),            //          .data
		.sink2_startofpacket (width_adapter_009_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket   (width_adapter_009_src_endofpacket),     //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (width_adapter_007_src_ready),           //     sink1.ready
		.sink1_valid          (width_adapter_007_src_valid),           //          .valid
		.sink1_channel        (width_adapter_007_src_channel),         //          .channel
		.sink1_data           (width_adapter_007_src_data),            //          .data
		.sink1_startofpacket  (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket    (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink2_ready          (width_adapter_010_src_ready),           //     sink2.ready
		.sink2_valid          (width_adapter_010_src_valid),           //          .valid
		.sink2_channel        (width_adapter_010_src_channel),         //          .channel
		.sink2_data           (width_adapter_010_src_data),            //          .data
		.sink2_startofpacket  (width_adapter_010_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket    (width_adapter_010_src_endofpacket),     //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src1_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src1_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (crosser_001_out_ready),                 //     sink6.ready
		.sink6_valid          (crosser_001_out_valid),                 //          .valid
		.sink6_channel        (crosser_001_out_channel),               //          .channel
		.sink6_data           (crosser_001_out_data),                  //          .data
		.sink6_startofpacket  (crosser_001_out_startofpacket),         //          .startofpacket
		.sink6_endofpacket    (crosser_001_out_endofpacket),           //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (rsp_xbar_demux_015_src0_ready),         //    sink15.ready
		.sink15_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink15_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink15_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.sink15_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink15_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios2_rsp_xbar_mux rsp_xbar_mux_002 (
		.clk                 (altpll_c0_clk),                         //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_008_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_008_src_valid),           //          .valid
		.sink0_channel       (width_adapter_008_src_channel),         //          .channel
		.sink0_data          (width_adapter_008_src_data),            //          .data
		.sink0_startofpacket (width_adapter_008_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_008_src_endofpacket),     //          .endofpacket
		.sink1_ready         (width_adapter_011_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_011_src_valid),           //          .valid
		.sink1_channel       (width_adapter_011_src_channel),         //          .channel
		.sink1_data          (width_adapter_011_src_data),            //          .data
		.sink1_startofpacket (width_adapter_011_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_011_src_endofpacket),     //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_010_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_015_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_015_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_015_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_015_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_015_src1_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (altpll_c0_clk),                     //       clk.clk
		.reset                (rst_controller_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_src1_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_src_data),            //          .data
		.out_channel          (width_adapter_src_channel),         //          .channel
		.out_valid            (width_adapter_src_valid),           //          .valid
		.out_ready            (width_adapter_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                             // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_001 (
		.clk                  (altpll_c0_clk),                       //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src2_valid),           //      sink.valid
		.in_channel           (cmd_xbar_demux_src2_channel),         //          .channel
		.in_startofpacket     (cmd_xbar_demux_src2_startofpacket),   //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src2_endofpacket),     //          .endofpacket
		.in_ready             (cmd_xbar_demux_src2_ready),           //          .ready
		.in_data              (cmd_xbar_demux_src2_data),            //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src1_data),          //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_002_src_data),            //          .data
		.out_channel          (width_adapter_002_src_channel),         //          .channel
		.out_valid            (width_adapter_002_src_valid),           //          .valid
		.out_ready            (width_adapter_002_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_003 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src2_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src2_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src2_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src2_data),          //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_003_src_data),            //          .data
		.out_channel          (width_adapter_003_src_channel),         //          .channel
		.out_valid            (width_adapter_003_src_valid),           //          .valid
		.out_ready            (width_adapter_003_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_004 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_002_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_004_src_data),            //          .data
		.out_channel          (width_adapter_004_src_channel),         //          .channel
		.out_valid            (width_adapter_004_src_valid),           //          .valid
		.out_ready            (width_adapter_004_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (88),
		.OUT_PKT_RESPONSE_STATUS_L     (87),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (89),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_005 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_002_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_002_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_002_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_002_src1_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_006 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_001_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_001_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_001_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_001_src0_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_006_src_data),            //          .data
		.out_channel          (width_adapter_006_src_channel),         //          .channel
		.out_valid            (width_adapter_006_src_valid),           //          .valid
		.out_ready            (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_007 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_001_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_001_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_001_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_001_src1_data),          //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_007_src_data),            //          .data
		.out_channel          (width_adapter_007_src_channel),         //          .channel
		.out_valid            (width_adapter_007_src_valid),           //          .valid
		.out_ready            (width_adapter_007_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_008 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_001_src2_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_001_src2_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_001_src2_ready),         //          .ready
		.in_data              (rsp_xbar_demux_001_src2_data),          //          .data
		.out_endofpacket      (width_adapter_008_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_008_src_data),            //          .data
		.out_channel          (width_adapter_008_src_channel),         //          .channel
		.out_valid            (width_adapter_008_src_valid),           //          .valid
		.out_ready            (width_adapter_008_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_008_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_009 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src0_data),          //          .data
		.out_endofpacket      (width_adapter_009_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_009_src_data),            //          .data
		.out_channel          (width_adapter_009_src_channel),         //          .channel
		.out_valid            (width_adapter_009_src_valid),           //          .valid
		.out_ready            (width_adapter_009_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_009_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_010 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src1_data),          //          .data
		.out_endofpacket      (width_adapter_010_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_010_src_data),            //          .data
		.out_channel          (width_adapter_010_src_channel),         //          .channel
		.out_valid            (width_adapter_010_src_valid),           //          .valid
		.out_ready            (width_adapter_010_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_010_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (88),
		.IN_PKT_RESPONSE_STATUS_L      (87),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (89),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (16),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_011 (
		.clk                  (altpll_c0_clk),                         //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_002_src2_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_002_src2_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_002_src2_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_002_src2_ready),         //          .ready
		.in_data              (rsp_xbar_demux_002_src2_data),          //          .data
		.out_endofpacket      (width_adapter_011_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_011_src_data),            //          .data
		.out_channel          (width_adapter_011_src_channel),         //          .channel
		.out_valid            (width_adapter_011_src_valid),           //          .valid
		.out_ready            (width_adapter_011_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_011_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (altpll_c0_clk),                         //        in_clk.clk
		.in_reset          (rst_controller_reset_out_reset),        //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src6_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src6_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src6_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src6_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src6_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (16),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (altpll_c0_clk),                         //       out_clk.clk
		.out_reset         (rst_controller_reset_out_reset),        // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_006_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_006_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_006_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_006_src0_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	nios2_irq_mapper irq_mapper (
		.clk           (altpll_c0_clk),                  //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),       // receiver8.irq
		.receiver9_irq (irq_mapper_receiver9_irq),       // receiver9.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

endmodule
